/home/linux/ieng6/ee260bwi25/sparanjpay/ECE260B_Project/dual_core/pnr/core/subckt/sram_w8_64b.lef