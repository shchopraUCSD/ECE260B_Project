##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 00:57:38 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w8_160b
  CLASS BLOCK ;
  SIZE 181.2000 BY 180.4000 ;
  FOREIGN sram_w8_160b 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 78.3500 0.6000 78.4500 ;
    END
  END CLK
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.8500 0.0000 169.9500 0.6000 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 0.0000 168.9500 0.6000 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.8500 0.0000 167.9500 0.6000 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 0.0000 166.9500 0.6000 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.8500 0.0000 165.9500 0.6000 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 0.0000 164.9500 0.6000 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 0.0000 163.9500 0.6000 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 0.0000 162.9500 0.6000 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.8500 0.0000 161.9500 0.6000 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 0.0000 160.9500 0.6000 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.8500 0.0000 159.9500 0.6000 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 0.0000 158.9500 0.6000 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.8500 0.0000 157.9500 0.6000 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 0.0000 156.9500 0.6000 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 0.0000 155.9500 0.6000 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 0.0000 154.9500 0.6000 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.8500 0.0000 153.9500 0.6000 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 0.0000 152.9500 0.6000 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.8500 0.0000 151.9500 0.6000 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 0.0000 150.9500 0.6000 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.8500 0.0000 149.9500 0.6000 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 0.0000 148.9500 0.6000 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.8500 0.0000 147.9500 0.6000 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 0.0000 146.9500 0.6000 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.8500 0.0000 145.9500 0.6000 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 0.0000 144.9500 0.6000 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.8500 0.0000 143.9500 0.6000 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 0.0000 142.9500 0.6000 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.8500 0.0000 141.9500 0.6000 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 0.0000 140.9500 0.6000 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.8500 0.0000 139.9500 0.6000 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 0.0000 138.9500 0.6000 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.8500 0.0000 137.9500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 0.0000 136.9500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.8500 0.0000 135.9500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 0.0000 134.9500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.8500 0.0000 133.9500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 0.0000 132.9500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.8500 0.0000 131.9500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 0.0000 130.9500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.8500 0.0000 129.9500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 0.0000 128.9500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.8500 0.0000 127.9500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 0.0000 126.9500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.8500 0.0000 125.9500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 0.0000 124.9500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.8500 0.0000 123.9500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 0.0000 122.9500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.8500 0.0000 121.9500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.8500 0.0000 120.9500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.8500 0.0000 119.9500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 0.0000 118.9500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.8500 0.0000 117.9500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.8500 0.0000 116.9500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.8500 0.0000 115.9500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 0.0000 114.9500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.8500 0.0000 113.9500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.8500 0.0000 112.9500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.8500 0.0000 111.9500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 0.0000 110.9500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.8500 0.0000 109.9500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.8500 0.0000 108.9500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.8500 0.0000 107.9500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 0.0000 106.9500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.8500 0.0000 105.9500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.8500 0.0000 104.9500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.8500 0.0000 103.9500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 0.0000 102.9500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.8500 0.0000 101.9500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.8500 0.0000 100.9500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.8500 0.0000 99.9500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 0.0000 98.9500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.8500 0.0000 97.9500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.8500 0.0000 96.9500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.8500 0.0000 95.9500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 0.0000 94.9500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.8500 0.0000 93.9500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.8500 0.0000 92.9500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.8500 0.0000 91.9500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 0.0000 90.9500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.8500 0.0000 89.9500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.8500 0.0000 88.9500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.8500 0.0000 87.9500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 0.0000 86.9500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.8500 0.0000 85.9500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.8500 0.0000 84.9500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.8500 0.0000 83.9500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 0.0000 82.9500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.8500 0.0000 81.9500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.8500 0.0000 80.9500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.8500 0.0000 79.9500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 0.0000 78.9500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.8500 0.0000 77.9500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.8500 0.0000 76.9500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.8500 0.0000 75.9500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 0.0000 74.9500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.8500 0.0000 73.9500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.8500 0.0000 72.9500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.8500 0.0000 71.9500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 0.0000 70.9500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.8500 0.0000 69.9500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.8500 0.0000 68.9500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.8500 0.0000 67.9500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 0.0000 66.9500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.8500 0.0000 65.9500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.8500 0.0000 64.9500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.8500 0.0000 63.9500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 0.0000 62.9500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.8500 0.0000 61.9500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.8500 0.0000 60.9500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.8500 0.0000 59.9500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 0.0000 58.9500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.8500 0.0000 57.9500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.8500 0.0000 56.9500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.8500 0.0000 55.9500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 0.0000 54.9500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.8500 0.0000 53.9500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.8500 0.0000 52.9500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.8500 0.0000 51.9500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 0.0000 50.9500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.8500 0.0000 49.9500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.8500 0.0000 48.9500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.8500 0.0000 47.9500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 0.0000 46.9500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.8500 0.0000 45.9500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.8500 0.0000 44.9500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.8500 0.0000 43.9500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 0.0000 42.9500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.8500 0.0000 41.9500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 0.0000 40.9500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.8500 0.0000 39.9500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 0.0000 38.9500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.8500 0.0000 37.9500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8500 0.0000 36.9500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.8500 0.0000 35.9500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 0.0000 34.9500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.8500 0.0000 33.9500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.8500 0.0000 32.9500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.8500 0.0000 31.9500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 0.0000 30.9500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8500 0.0000 29.9500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8500 0.0000 28.9500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.8500 0.0000 27.9500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 0.0000 26.9500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8500 0.0000 25.9500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8500 0.0000 24.9500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.8500 0.0000 23.9500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 0.0000 22.9500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.8500 0.0000 21.9500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8500 0.0000 20.9500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8500 0.0000 19.9500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 0.0000 18.9500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.8500 0.0000 17.9500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8500 0.0000 16.9500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.8500 0.0000 15.9500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.8500 0.0000 14.9500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.8500 0.0000 13.9500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.8500 0.0000 12.9500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.8500 0.0000 11.9500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.8500 0.0000 10.9500 0.6000 ;
    END
  END D[0]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.8500 179.8000 169.9500 180.4000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 179.8000 168.9500 180.4000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.8500 179.8000 167.9500 180.4000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 179.8000 166.9500 180.4000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.8500 179.8000 165.9500 180.4000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 179.8000 164.9500 180.4000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 179.8000 163.9500 180.4000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 179.8000 162.9500 180.4000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.8500 179.8000 161.9500 180.4000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 179.8000 160.9500 180.4000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.8500 179.8000 159.9500 180.4000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 179.8000 158.9500 180.4000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.8500 179.8000 157.9500 180.4000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 179.8000 156.9500 180.4000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 179.8000 155.9500 180.4000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 179.8000 154.9500 180.4000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.8500 179.8000 153.9500 180.4000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 179.8000 152.9500 180.4000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.8500 179.8000 151.9500 180.4000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 179.8000 150.9500 180.4000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.8500 179.8000 149.9500 180.4000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 179.8000 148.9500 180.4000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.8500 179.8000 147.9500 180.4000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 179.8000 146.9500 180.4000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.8500 179.8000 145.9500 180.4000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 179.8000 144.9500 180.4000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.8500 179.8000 143.9500 180.4000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 179.8000 142.9500 180.4000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.8500 179.8000 141.9500 180.4000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 179.8000 140.9500 180.4000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.8500 179.8000 139.9500 180.4000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 179.8000 138.9500 180.4000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.8500 179.8000 137.9500 180.4000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 179.8000 136.9500 180.4000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.8500 179.8000 135.9500 180.4000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 179.8000 134.9500 180.4000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.8500 179.8000 133.9500 180.4000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 179.8000 132.9500 180.4000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.8500 179.8000 131.9500 180.4000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 179.8000 130.9500 180.4000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.8500 179.8000 129.9500 180.4000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 179.8000 128.9500 180.4000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.8500 179.8000 127.9500 180.4000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 179.8000 126.9500 180.4000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.8500 179.8000 125.9500 180.4000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 179.8000 124.9500 180.4000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.8500 179.8000 123.9500 180.4000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 179.8000 122.9500 180.4000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.8500 179.8000 121.9500 180.4000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.8500 179.8000 120.9500 180.4000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.8500 179.8000 119.9500 180.4000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 179.8000 118.9500 180.4000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.8500 179.8000 117.9500 180.4000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.8500 179.8000 116.9500 180.4000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.8500 179.8000 115.9500 180.4000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 179.8000 114.9500 180.4000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.8500 179.8000 113.9500 180.4000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.8500 179.8000 112.9500 180.4000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.8500 179.8000 111.9500 180.4000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 179.8000 110.9500 180.4000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.8500 179.8000 109.9500 180.4000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.8500 179.8000 108.9500 180.4000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.8500 179.8000 107.9500 180.4000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 179.8000 106.9500 180.4000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.8500 179.8000 105.9500 180.4000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.8500 179.8000 104.9500 180.4000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.8500 179.8000 103.9500 180.4000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 179.8000 102.9500 180.4000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.8500 179.8000 101.9500 180.4000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.8500 179.8000 100.9500 180.4000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.8500 179.8000 99.9500 180.4000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 179.8000 98.9500 180.4000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.8500 179.8000 97.9500 180.4000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.8500 179.8000 96.9500 180.4000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.8500 179.8000 95.9500 180.4000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 179.8000 94.9500 180.4000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.8500 179.8000 93.9500 180.4000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.8500 179.8000 92.9500 180.4000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.8500 179.8000 91.9500 180.4000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 179.8000 90.9500 180.4000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.8500 179.8000 89.9500 180.4000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.8500 179.8000 88.9500 180.4000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.8500 179.8000 87.9500 180.4000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.8500 179.8000 86.9500 180.4000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.8500 179.8000 85.9500 180.4000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.8500 179.8000 84.9500 180.4000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.8500 179.8000 83.9500 180.4000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.8500 179.8000 82.9500 180.4000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.8500 179.8000 81.9500 180.4000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.8500 179.8000 80.9500 180.4000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.8500 179.8000 79.9500 180.4000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.8500 179.8000 78.9500 180.4000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.8500 179.8000 77.9500 180.4000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.8500 179.8000 76.9500 180.4000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.8500 179.8000 75.9500 180.4000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.8500 179.8000 74.9500 180.4000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.8500 179.8000 73.9500 180.4000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.8500 179.8000 72.9500 180.4000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.8500 179.8000 71.9500 180.4000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.8500 179.8000 70.9500 180.4000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.8500 179.8000 69.9500 180.4000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.8500 179.8000 68.9500 180.4000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.8500 179.8000 67.9500 180.4000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.8500 179.8000 66.9500 180.4000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.8500 179.8000 65.9500 180.4000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.8500 179.8000 64.9500 180.4000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.8500 179.8000 63.9500 180.4000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.8500 179.8000 62.9500 180.4000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.8500 179.8000 61.9500 180.4000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.8500 179.8000 60.9500 180.4000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.8500 179.8000 59.9500 180.4000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.8500 179.8000 58.9500 180.4000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.8500 179.8000 57.9500 180.4000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.8500 179.8000 56.9500 180.4000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.8500 179.8000 55.9500 180.4000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.8500 179.8000 54.9500 180.4000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.8500 179.8000 53.9500 180.4000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.8500 179.8000 52.9500 180.4000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.8500 179.8000 51.9500 180.4000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.8500 179.8000 50.9500 180.4000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.8500 179.8000 49.9500 180.4000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.8500 179.8000 48.9500 180.4000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.8500 179.8000 47.9500 180.4000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.8500 179.8000 46.9500 180.4000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.8500 179.8000 45.9500 180.4000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.8500 179.8000 44.9500 180.4000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.8500 179.8000 43.9500 180.4000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.8500 179.8000 42.9500 180.4000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.8500 179.8000 41.9500 180.4000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 179.8000 40.9500 180.4000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.8500 179.8000 39.9500 180.4000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.8500 179.8000 38.9500 180.4000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.8500 179.8000 37.9500 180.4000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.8500 179.8000 36.9500 180.4000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.8500 179.8000 35.9500 180.4000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.8500 179.8000 34.9500 180.4000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.8500 179.8000 33.9500 180.4000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.8500 179.8000 32.9500 180.4000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.8500 179.8000 31.9500 180.4000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.8500 179.8000 30.9500 180.4000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.8500 179.8000 29.9500 180.4000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.8500 179.8000 28.9500 180.4000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.8500 179.8000 27.9500 180.4000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.8500 179.8000 26.9500 180.4000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.8500 179.8000 25.9500 180.4000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.8500 179.8000 24.9500 180.4000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.8500 179.8000 23.9500 180.4000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.8500 179.8000 22.9500 180.4000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.8500 179.8000 21.9500 180.4000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.8500 179.8000 20.9500 180.4000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8500 179.8000 19.9500 180.4000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.8500 179.8000 18.9500 180.4000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.8500 179.8000 17.9500 180.4000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.8500 179.8000 16.9500 180.4000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.8500 179.8000 15.9500 180.4000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.8500 179.8000 14.9500 180.4000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.8500 179.8000 13.9500 180.4000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.8500 179.8000 12.9500 180.4000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.8500 179.8000 11.9500 180.4000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.8500 179.8000 10.9500 180.4000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 86.3500 0.6000 86.4500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 82.3500 0.6000 82.4500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 90.3500 0.6000 90.4500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 94.3500 0.6000 94.4500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 98.3500 0.6000 98.4500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 102.3500 0.6000 102.4500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 44.4400 2.0000 46.4400 178.4000 ;
        RECT 28.2200 2.0000 30.2200 178.4000 ;
        RECT 12.0000 2.0000 14.0000 178.4000 ;
        RECT 76.8800 2.0000 78.8800 178.4000 ;
        RECT 60.6600 2.0000 62.6600 178.4000 ;
        RECT 125.5400 2.0000 127.5400 178.4000 ;
        RECT 109.3200 2.0000 111.3200 178.4000 ;
        RECT 93.1000 2.0000 95.1000 178.4000 ;
        RECT 157.9800 2.0000 159.9800 178.4000 ;
        RECT 141.7600 2.0000 143.7600 178.4000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 37.4400 2.0000 39.4400 178.4000 ;
        RECT 21.2200 2.0000 23.2200 178.4000 ;
        RECT 5.0000 2.0000 7.0000 178.4000 ;
        RECT 86.1000 2.0000 88.1000 178.4000 ;
        RECT 69.8800 2.0000 71.8800 178.4000 ;
        RECT 53.6600 2.0000 55.6600 178.4000 ;
        RECT 134.7600 2.0000 136.7600 178.4000 ;
        RECT 118.5400 2.0000 120.5400 178.4000 ;
        RECT 102.3200 2.0000 104.3200 178.4000 ;
        RECT 150.9800 2.0000 152.9800 178.4000 ;
        RECT 21.2200 1.8350 23.2200 2.1650 ;
        RECT 5.0000 1.8350 7.0000 2.1650 ;
        RECT 37.4400 1.8350 39.4400 2.1650 ;
        RECT 53.6600 1.8350 55.6600 2.1650 ;
        RECT 69.8800 1.8350 71.8800 2.1650 ;
        RECT 86.1000 1.8350 88.1000 2.1650 ;
        RECT 134.7600 1.8350 136.7600 2.1650 ;
        RECT 102.3200 1.8350 104.3200 2.1650 ;
        RECT 118.5400 1.8350 120.5400 2.1650 ;
        RECT 150.9800 1.8350 152.9800 2.1650 ;
        RECT 21.2200 178.2350 23.2200 178.5650 ;
        RECT 5.0000 178.2350 7.0000 178.5650 ;
        RECT 37.4400 178.2350 39.4400 178.5650 ;
        RECT 53.6600 178.2350 55.6600 178.5650 ;
        RECT 69.8800 178.2350 71.8800 178.5650 ;
        RECT 86.1000 178.2350 88.1000 178.5650 ;
        RECT 134.7600 178.2350 136.7600 178.5650 ;
        RECT 102.3200 178.2350 104.3200 178.5650 ;
        RECT 118.5400 178.2350 120.5400 178.5650 ;
        RECT 150.9800 178.2350 152.9800 178.5650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 181.2000 180.4000 ;
    LAYER M2 ;
      RECT 170.0500 179.7000 181.2000 180.4000 ;
      RECT 169.0500 179.7000 169.7500 180.4000 ;
      RECT 168.0500 179.7000 168.7500 180.4000 ;
      RECT 167.0500 179.7000 167.7500 180.4000 ;
      RECT 166.0500 179.7000 166.7500 180.4000 ;
      RECT 165.0500 179.7000 165.7500 180.4000 ;
      RECT 164.0500 179.7000 164.7500 180.4000 ;
      RECT 163.0500 179.7000 163.7500 180.4000 ;
      RECT 162.0500 179.7000 162.7500 180.4000 ;
      RECT 161.0500 179.7000 161.7500 180.4000 ;
      RECT 160.0500 179.7000 160.7500 180.4000 ;
      RECT 159.0500 179.7000 159.7500 180.4000 ;
      RECT 158.0500 179.7000 158.7500 180.4000 ;
      RECT 157.0500 179.7000 157.7500 180.4000 ;
      RECT 156.0500 179.7000 156.7500 180.4000 ;
      RECT 155.0500 179.7000 155.7500 180.4000 ;
      RECT 154.0500 179.7000 154.7500 180.4000 ;
      RECT 153.0500 179.7000 153.7500 180.4000 ;
      RECT 152.0500 179.7000 152.7500 180.4000 ;
      RECT 151.0500 179.7000 151.7500 180.4000 ;
      RECT 150.0500 179.7000 150.7500 180.4000 ;
      RECT 149.0500 179.7000 149.7500 180.4000 ;
      RECT 148.0500 179.7000 148.7500 180.4000 ;
      RECT 147.0500 179.7000 147.7500 180.4000 ;
      RECT 146.0500 179.7000 146.7500 180.4000 ;
      RECT 145.0500 179.7000 145.7500 180.4000 ;
      RECT 144.0500 179.7000 144.7500 180.4000 ;
      RECT 143.0500 179.7000 143.7500 180.4000 ;
      RECT 142.0500 179.7000 142.7500 180.4000 ;
      RECT 141.0500 179.7000 141.7500 180.4000 ;
      RECT 140.0500 179.7000 140.7500 180.4000 ;
      RECT 139.0500 179.7000 139.7500 180.4000 ;
      RECT 138.0500 179.7000 138.7500 180.4000 ;
      RECT 137.0500 179.7000 137.7500 180.4000 ;
      RECT 136.0500 179.7000 136.7500 180.4000 ;
      RECT 135.0500 179.7000 135.7500 180.4000 ;
      RECT 134.0500 179.7000 134.7500 180.4000 ;
      RECT 133.0500 179.7000 133.7500 180.4000 ;
      RECT 132.0500 179.7000 132.7500 180.4000 ;
      RECT 131.0500 179.7000 131.7500 180.4000 ;
      RECT 130.0500 179.7000 130.7500 180.4000 ;
      RECT 129.0500 179.7000 129.7500 180.4000 ;
      RECT 128.0500 179.7000 128.7500 180.4000 ;
      RECT 127.0500 179.7000 127.7500 180.4000 ;
      RECT 126.0500 179.7000 126.7500 180.4000 ;
      RECT 125.0500 179.7000 125.7500 180.4000 ;
      RECT 124.0500 179.7000 124.7500 180.4000 ;
      RECT 123.0500 179.7000 123.7500 180.4000 ;
      RECT 122.0500 179.7000 122.7500 180.4000 ;
      RECT 121.0500 179.7000 121.7500 180.4000 ;
      RECT 120.0500 179.7000 120.7500 180.4000 ;
      RECT 119.0500 179.7000 119.7500 180.4000 ;
      RECT 118.0500 179.7000 118.7500 180.4000 ;
      RECT 117.0500 179.7000 117.7500 180.4000 ;
      RECT 116.0500 179.7000 116.7500 180.4000 ;
      RECT 115.0500 179.7000 115.7500 180.4000 ;
      RECT 114.0500 179.7000 114.7500 180.4000 ;
      RECT 113.0500 179.7000 113.7500 180.4000 ;
      RECT 112.0500 179.7000 112.7500 180.4000 ;
      RECT 111.0500 179.7000 111.7500 180.4000 ;
      RECT 110.0500 179.7000 110.7500 180.4000 ;
      RECT 109.0500 179.7000 109.7500 180.4000 ;
      RECT 108.0500 179.7000 108.7500 180.4000 ;
      RECT 107.0500 179.7000 107.7500 180.4000 ;
      RECT 106.0500 179.7000 106.7500 180.4000 ;
      RECT 105.0500 179.7000 105.7500 180.4000 ;
      RECT 104.0500 179.7000 104.7500 180.4000 ;
      RECT 103.0500 179.7000 103.7500 180.4000 ;
      RECT 102.0500 179.7000 102.7500 180.4000 ;
      RECT 101.0500 179.7000 101.7500 180.4000 ;
      RECT 100.0500 179.7000 100.7500 180.4000 ;
      RECT 99.0500 179.7000 99.7500 180.4000 ;
      RECT 98.0500 179.7000 98.7500 180.4000 ;
      RECT 97.0500 179.7000 97.7500 180.4000 ;
      RECT 96.0500 179.7000 96.7500 180.4000 ;
      RECT 95.0500 179.7000 95.7500 180.4000 ;
      RECT 94.0500 179.7000 94.7500 180.4000 ;
      RECT 93.0500 179.7000 93.7500 180.4000 ;
      RECT 92.0500 179.7000 92.7500 180.4000 ;
      RECT 91.0500 179.7000 91.7500 180.4000 ;
      RECT 90.0500 179.7000 90.7500 180.4000 ;
      RECT 89.0500 179.7000 89.7500 180.4000 ;
      RECT 88.0500 179.7000 88.7500 180.4000 ;
      RECT 87.0500 179.7000 87.7500 180.4000 ;
      RECT 86.0500 179.7000 86.7500 180.4000 ;
      RECT 85.0500 179.7000 85.7500 180.4000 ;
      RECT 84.0500 179.7000 84.7500 180.4000 ;
      RECT 83.0500 179.7000 83.7500 180.4000 ;
      RECT 82.0500 179.7000 82.7500 180.4000 ;
      RECT 81.0500 179.7000 81.7500 180.4000 ;
      RECT 80.0500 179.7000 80.7500 180.4000 ;
      RECT 79.0500 179.7000 79.7500 180.4000 ;
      RECT 78.0500 179.7000 78.7500 180.4000 ;
      RECT 77.0500 179.7000 77.7500 180.4000 ;
      RECT 76.0500 179.7000 76.7500 180.4000 ;
      RECT 75.0500 179.7000 75.7500 180.4000 ;
      RECT 74.0500 179.7000 74.7500 180.4000 ;
      RECT 73.0500 179.7000 73.7500 180.4000 ;
      RECT 72.0500 179.7000 72.7500 180.4000 ;
      RECT 71.0500 179.7000 71.7500 180.4000 ;
      RECT 70.0500 179.7000 70.7500 180.4000 ;
      RECT 69.0500 179.7000 69.7500 180.4000 ;
      RECT 68.0500 179.7000 68.7500 180.4000 ;
      RECT 67.0500 179.7000 67.7500 180.4000 ;
      RECT 66.0500 179.7000 66.7500 180.4000 ;
      RECT 65.0500 179.7000 65.7500 180.4000 ;
      RECT 64.0500 179.7000 64.7500 180.4000 ;
      RECT 63.0500 179.7000 63.7500 180.4000 ;
      RECT 62.0500 179.7000 62.7500 180.4000 ;
      RECT 61.0500 179.7000 61.7500 180.4000 ;
      RECT 60.0500 179.7000 60.7500 180.4000 ;
      RECT 59.0500 179.7000 59.7500 180.4000 ;
      RECT 58.0500 179.7000 58.7500 180.4000 ;
      RECT 57.0500 179.7000 57.7500 180.4000 ;
      RECT 56.0500 179.7000 56.7500 180.4000 ;
      RECT 55.0500 179.7000 55.7500 180.4000 ;
      RECT 54.0500 179.7000 54.7500 180.4000 ;
      RECT 53.0500 179.7000 53.7500 180.4000 ;
      RECT 52.0500 179.7000 52.7500 180.4000 ;
      RECT 51.0500 179.7000 51.7500 180.4000 ;
      RECT 50.0500 179.7000 50.7500 180.4000 ;
      RECT 49.0500 179.7000 49.7500 180.4000 ;
      RECT 48.0500 179.7000 48.7500 180.4000 ;
      RECT 47.0500 179.7000 47.7500 180.4000 ;
      RECT 46.0500 179.7000 46.7500 180.4000 ;
      RECT 45.0500 179.7000 45.7500 180.4000 ;
      RECT 44.0500 179.7000 44.7500 180.4000 ;
      RECT 43.0500 179.7000 43.7500 180.4000 ;
      RECT 42.0500 179.7000 42.7500 180.4000 ;
      RECT 41.0500 179.7000 41.7500 180.4000 ;
      RECT 40.0500 179.7000 40.7500 180.4000 ;
      RECT 39.0500 179.7000 39.7500 180.4000 ;
      RECT 38.0500 179.7000 38.7500 180.4000 ;
      RECT 37.0500 179.7000 37.7500 180.4000 ;
      RECT 36.0500 179.7000 36.7500 180.4000 ;
      RECT 35.0500 179.7000 35.7500 180.4000 ;
      RECT 34.0500 179.7000 34.7500 180.4000 ;
      RECT 33.0500 179.7000 33.7500 180.4000 ;
      RECT 32.0500 179.7000 32.7500 180.4000 ;
      RECT 31.0500 179.7000 31.7500 180.4000 ;
      RECT 30.0500 179.7000 30.7500 180.4000 ;
      RECT 29.0500 179.7000 29.7500 180.4000 ;
      RECT 28.0500 179.7000 28.7500 180.4000 ;
      RECT 27.0500 179.7000 27.7500 180.4000 ;
      RECT 26.0500 179.7000 26.7500 180.4000 ;
      RECT 25.0500 179.7000 25.7500 180.4000 ;
      RECT 24.0500 179.7000 24.7500 180.4000 ;
      RECT 23.0500 179.7000 23.7500 180.4000 ;
      RECT 22.0500 179.7000 22.7500 180.4000 ;
      RECT 21.0500 179.7000 21.7500 180.4000 ;
      RECT 20.0500 179.7000 20.7500 180.4000 ;
      RECT 19.0500 179.7000 19.7500 180.4000 ;
      RECT 18.0500 179.7000 18.7500 180.4000 ;
      RECT 17.0500 179.7000 17.7500 180.4000 ;
      RECT 16.0500 179.7000 16.7500 180.4000 ;
      RECT 15.0500 179.7000 15.7500 180.4000 ;
      RECT 14.0500 179.7000 14.7500 180.4000 ;
      RECT 13.0500 179.7000 13.7500 180.4000 ;
      RECT 12.0500 179.7000 12.7500 180.4000 ;
      RECT 11.0500 179.7000 11.7500 180.4000 ;
      RECT 0.0000 179.7000 10.7500 180.4000 ;
      RECT 0.0000 0.7000 181.2000 179.7000 ;
      RECT 170.0500 0.0000 181.2000 0.7000 ;
      RECT 169.0500 0.0000 169.7500 0.7000 ;
      RECT 168.0500 0.0000 168.7500 0.7000 ;
      RECT 167.0500 0.0000 167.7500 0.7000 ;
      RECT 166.0500 0.0000 166.7500 0.7000 ;
      RECT 165.0500 0.0000 165.7500 0.7000 ;
      RECT 164.0500 0.0000 164.7500 0.7000 ;
      RECT 163.0500 0.0000 163.7500 0.7000 ;
      RECT 162.0500 0.0000 162.7500 0.7000 ;
      RECT 161.0500 0.0000 161.7500 0.7000 ;
      RECT 160.0500 0.0000 160.7500 0.7000 ;
      RECT 159.0500 0.0000 159.7500 0.7000 ;
      RECT 158.0500 0.0000 158.7500 0.7000 ;
      RECT 157.0500 0.0000 157.7500 0.7000 ;
      RECT 156.0500 0.0000 156.7500 0.7000 ;
      RECT 155.0500 0.0000 155.7500 0.7000 ;
      RECT 154.0500 0.0000 154.7500 0.7000 ;
      RECT 153.0500 0.0000 153.7500 0.7000 ;
      RECT 152.0500 0.0000 152.7500 0.7000 ;
      RECT 151.0500 0.0000 151.7500 0.7000 ;
      RECT 150.0500 0.0000 150.7500 0.7000 ;
      RECT 149.0500 0.0000 149.7500 0.7000 ;
      RECT 148.0500 0.0000 148.7500 0.7000 ;
      RECT 147.0500 0.0000 147.7500 0.7000 ;
      RECT 146.0500 0.0000 146.7500 0.7000 ;
      RECT 145.0500 0.0000 145.7500 0.7000 ;
      RECT 144.0500 0.0000 144.7500 0.7000 ;
      RECT 143.0500 0.0000 143.7500 0.7000 ;
      RECT 142.0500 0.0000 142.7500 0.7000 ;
      RECT 141.0500 0.0000 141.7500 0.7000 ;
      RECT 140.0500 0.0000 140.7500 0.7000 ;
      RECT 139.0500 0.0000 139.7500 0.7000 ;
      RECT 138.0500 0.0000 138.7500 0.7000 ;
      RECT 137.0500 0.0000 137.7500 0.7000 ;
      RECT 136.0500 0.0000 136.7500 0.7000 ;
      RECT 135.0500 0.0000 135.7500 0.7000 ;
      RECT 134.0500 0.0000 134.7500 0.7000 ;
      RECT 133.0500 0.0000 133.7500 0.7000 ;
      RECT 132.0500 0.0000 132.7500 0.7000 ;
      RECT 131.0500 0.0000 131.7500 0.7000 ;
      RECT 130.0500 0.0000 130.7500 0.7000 ;
      RECT 129.0500 0.0000 129.7500 0.7000 ;
      RECT 128.0500 0.0000 128.7500 0.7000 ;
      RECT 127.0500 0.0000 127.7500 0.7000 ;
      RECT 126.0500 0.0000 126.7500 0.7000 ;
      RECT 125.0500 0.0000 125.7500 0.7000 ;
      RECT 124.0500 0.0000 124.7500 0.7000 ;
      RECT 123.0500 0.0000 123.7500 0.7000 ;
      RECT 122.0500 0.0000 122.7500 0.7000 ;
      RECT 121.0500 0.0000 121.7500 0.7000 ;
      RECT 120.0500 0.0000 120.7500 0.7000 ;
      RECT 119.0500 0.0000 119.7500 0.7000 ;
      RECT 118.0500 0.0000 118.7500 0.7000 ;
      RECT 117.0500 0.0000 117.7500 0.7000 ;
      RECT 116.0500 0.0000 116.7500 0.7000 ;
      RECT 115.0500 0.0000 115.7500 0.7000 ;
      RECT 114.0500 0.0000 114.7500 0.7000 ;
      RECT 113.0500 0.0000 113.7500 0.7000 ;
      RECT 112.0500 0.0000 112.7500 0.7000 ;
      RECT 111.0500 0.0000 111.7500 0.7000 ;
      RECT 110.0500 0.0000 110.7500 0.7000 ;
      RECT 109.0500 0.0000 109.7500 0.7000 ;
      RECT 108.0500 0.0000 108.7500 0.7000 ;
      RECT 107.0500 0.0000 107.7500 0.7000 ;
      RECT 106.0500 0.0000 106.7500 0.7000 ;
      RECT 105.0500 0.0000 105.7500 0.7000 ;
      RECT 104.0500 0.0000 104.7500 0.7000 ;
      RECT 103.0500 0.0000 103.7500 0.7000 ;
      RECT 102.0500 0.0000 102.7500 0.7000 ;
      RECT 101.0500 0.0000 101.7500 0.7000 ;
      RECT 100.0500 0.0000 100.7500 0.7000 ;
      RECT 99.0500 0.0000 99.7500 0.7000 ;
      RECT 98.0500 0.0000 98.7500 0.7000 ;
      RECT 97.0500 0.0000 97.7500 0.7000 ;
      RECT 96.0500 0.0000 96.7500 0.7000 ;
      RECT 95.0500 0.0000 95.7500 0.7000 ;
      RECT 94.0500 0.0000 94.7500 0.7000 ;
      RECT 93.0500 0.0000 93.7500 0.7000 ;
      RECT 92.0500 0.0000 92.7500 0.7000 ;
      RECT 91.0500 0.0000 91.7500 0.7000 ;
      RECT 90.0500 0.0000 90.7500 0.7000 ;
      RECT 89.0500 0.0000 89.7500 0.7000 ;
      RECT 88.0500 0.0000 88.7500 0.7000 ;
      RECT 87.0500 0.0000 87.7500 0.7000 ;
      RECT 86.0500 0.0000 86.7500 0.7000 ;
      RECT 85.0500 0.0000 85.7500 0.7000 ;
      RECT 84.0500 0.0000 84.7500 0.7000 ;
      RECT 83.0500 0.0000 83.7500 0.7000 ;
      RECT 82.0500 0.0000 82.7500 0.7000 ;
      RECT 81.0500 0.0000 81.7500 0.7000 ;
      RECT 80.0500 0.0000 80.7500 0.7000 ;
      RECT 79.0500 0.0000 79.7500 0.7000 ;
      RECT 78.0500 0.0000 78.7500 0.7000 ;
      RECT 77.0500 0.0000 77.7500 0.7000 ;
      RECT 76.0500 0.0000 76.7500 0.7000 ;
      RECT 75.0500 0.0000 75.7500 0.7000 ;
      RECT 74.0500 0.0000 74.7500 0.7000 ;
      RECT 73.0500 0.0000 73.7500 0.7000 ;
      RECT 72.0500 0.0000 72.7500 0.7000 ;
      RECT 71.0500 0.0000 71.7500 0.7000 ;
      RECT 70.0500 0.0000 70.7500 0.7000 ;
      RECT 69.0500 0.0000 69.7500 0.7000 ;
      RECT 68.0500 0.0000 68.7500 0.7000 ;
      RECT 67.0500 0.0000 67.7500 0.7000 ;
      RECT 66.0500 0.0000 66.7500 0.7000 ;
      RECT 65.0500 0.0000 65.7500 0.7000 ;
      RECT 64.0500 0.0000 64.7500 0.7000 ;
      RECT 63.0500 0.0000 63.7500 0.7000 ;
      RECT 62.0500 0.0000 62.7500 0.7000 ;
      RECT 61.0500 0.0000 61.7500 0.7000 ;
      RECT 60.0500 0.0000 60.7500 0.7000 ;
      RECT 59.0500 0.0000 59.7500 0.7000 ;
      RECT 58.0500 0.0000 58.7500 0.7000 ;
      RECT 57.0500 0.0000 57.7500 0.7000 ;
      RECT 56.0500 0.0000 56.7500 0.7000 ;
      RECT 55.0500 0.0000 55.7500 0.7000 ;
      RECT 54.0500 0.0000 54.7500 0.7000 ;
      RECT 53.0500 0.0000 53.7500 0.7000 ;
      RECT 52.0500 0.0000 52.7500 0.7000 ;
      RECT 51.0500 0.0000 51.7500 0.7000 ;
      RECT 50.0500 0.0000 50.7500 0.7000 ;
      RECT 49.0500 0.0000 49.7500 0.7000 ;
      RECT 48.0500 0.0000 48.7500 0.7000 ;
      RECT 47.0500 0.0000 47.7500 0.7000 ;
      RECT 46.0500 0.0000 46.7500 0.7000 ;
      RECT 45.0500 0.0000 45.7500 0.7000 ;
      RECT 44.0500 0.0000 44.7500 0.7000 ;
      RECT 43.0500 0.0000 43.7500 0.7000 ;
      RECT 42.0500 0.0000 42.7500 0.7000 ;
      RECT 41.0500 0.0000 41.7500 0.7000 ;
      RECT 40.0500 0.0000 40.7500 0.7000 ;
      RECT 39.0500 0.0000 39.7500 0.7000 ;
      RECT 38.0500 0.0000 38.7500 0.7000 ;
      RECT 37.0500 0.0000 37.7500 0.7000 ;
      RECT 36.0500 0.0000 36.7500 0.7000 ;
      RECT 35.0500 0.0000 35.7500 0.7000 ;
      RECT 34.0500 0.0000 34.7500 0.7000 ;
      RECT 33.0500 0.0000 33.7500 0.7000 ;
      RECT 32.0500 0.0000 32.7500 0.7000 ;
      RECT 31.0500 0.0000 31.7500 0.7000 ;
      RECT 30.0500 0.0000 30.7500 0.7000 ;
      RECT 29.0500 0.0000 29.7500 0.7000 ;
      RECT 28.0500 0.0000 28.7500 0.7000 ;
      RECT 27.0500 0.0000 27.7500 0.7000 ;
      RECT 26.0500 0.0000 26.7500 0.7000 ;
      RECT 25.0500 0.0000 25.7500 0.7000 ;
      RECT 24.0500 0.0000 24.7500 0.7000 ;
      RECT 23.0500 0.0000 23.7500 0.7000 ;
      RECT 22.0500 0.0000 22.7500 0.7000 ;
      RECT 21.0500 0.0000 21.7500 0.7000 ;
      RECT 20.0500 0.0000 20.7500 0.7000 ;
      RECT 19.0500 0.0000 19.7500 0.7000 ;
      RECT 18.0500 0.0000 18.7500 0.7000 ;
      RECT 17.0500 0.0000 17.7500 0.7000 ;
      RECT 16.0500 0.0000 16.7500 0.7000 ;
      RECT 15.0500 0.0000 15.7500 0.7000 ;
      RECT 14.0500 0.0000 14.7500 0.7000 ;
      RECT 13.0500 0.0000 13.7500 0.7000 ;
      RECT 12.0500 0.0000 12.7500 0.7000 ;
      RECT 11.0500 0.0000 11.7500 0.7000 ;
      RECT 0.0000 0.0000 10.7500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 102.5500 181.2000 180.4000 ;
      RECT 0.7000 102.2500 181.2000 102.5500 ;
      RECT 0.0000 98.5500 181.2000 102.2500 ;
      RECT 0.7000 98.2500 181.2000 98.5500 ;
      RECT 0.0000 94.5500 181.2000 98.2500 ;
      RECT 0.7000 94.2500 181.2000 94.5500 ;
      RECT 0.0000 90.5500 181.2000 94.2500 ;
      RECT 0.7000 90.2500 181.2000 90.5500 ;
      RECT 0.0000 86.5500 181.2000 90.2500 ;
      RECT 0.7000 86.2500 181.2000 86.5500 ;
      RECT 0.0000 82.5500 181.2000 86.2500 ;
      RECT 0.7000 82.2500 181.2000 82.5500 ;
      RECT 0.0000 78.5500 181.2000 82.2500 ;
      RECT 0.7000 78.2500 181.2000 78.5500 ;
      RECT 0.0000 0.0000 181.2000 78.2500 ;
    LAYER M4 ;
      RECT 0.0000 179.0650 181.2000 180.4000 ;
      RECT 153.4800 178.9000 181.2000 179.0650 ;
      RECT 137.2600 178.9000 150.4800 179.0650 ;
      RECT 121.0400 178.9000 134.2600 179.0650 ;
      RECT 104.8200 178.9000 118.0400 179.0650 ;
      RECT 88.6000 178.9000 101.8200 179.0650 ;
      RECT 72.3800 178.9000 85.6000 179.0650 ;
      RECT 56.1600 178.9000 69.3800 179.0650 ;
      RECT 39.9400 178.9000 53.1600 179.0650 ;
      RECT 23.7200 178.9000 36.9400 179.0650 ;
      RECT 7.5000 178.9000 20.7200 179.0650 ;
      RECT 160.4800 1.5000 181.2000 178.9000 ;
      RECT 153.4800 1.5000 157.4800 178.9000 ;
      RECT 144.2600 1.5000 150.4800 178.9000 ;
      RECT 137.2600 1.5000 141.2600 178.9000 ;
      RECT 128.0400 1.5000 134.2600 178.9000 ;
      RECT 121.0400 1.5000 125.0400 178.9000 ;
      RECT 111.8200 1.5000 118.0400 178.9000 ;
      RECT 104.8200 1.5000 108.8200 178.9000 ;
      RECT 95.6000 1.5000 101.8200 178.9000 ;
      RECT 88.6000 1.5000 92.6000 178.9000 ;
      RECT 79.3800 1.5000 85.6000 178.9000 ;
      RECT 72.3800 1.5000 76.3800 178.9000 ;
      RECT 63.1600 1.5000 69.3800 178.9000 ;
      RECT 56.1600 1.5000 60.1600 178.9000 ;
      RECT 46.9400 1.5000 53.1600 178.9000 ;
      RECT 39.9400 1.5000 43.9400 178.9000 ;
      RECT 30.7200 1.5000 36.9400 178.9000 ;
      RECT 23.7200 1.5000 27.7200 178.9000 ;
      RECT 14.5000 1.5000 20.7200 178.9000 ;
      RECT 7.5000 1.5000 11.5000 178.9000 ;
      RECT 153.4800 1.3350 181.2000 1.5000 ;
      RECT 137.2600 1.3350 150.4800 1.5000 ;
      RECT 121.0400 1.3350 134.2600 1.5000 ;
      RECT 104.8200 1.3350 118.0400 1.5000 ;
      RECT 88.6000 1.3350 101.8200 1.5000 ;
      RECT 72.3800 1.3350 85.6000 1.5000 ;
      RECT 56.1600 1.3350 69.3800 1.5000 ;
      RECT 39.9400 1.3350 53.1600 1.5000 ;
      RECT 23.7200 1.3350 36.9400 1.5000 ;
      RECT 7.5000 1.3350 20.7200 1.5000 ;
      RECT 0.0000 1.3350 4.5000 179.0650 ;
      RECT 0.0000 0.0000 181.2000 1.3350 ;
  END
END sram_w8_160b

END LIBRARY
