##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Wed Mar 19 19:53:11 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 639.8000 BY 639.2000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 325.3500 0.5200 325.4500 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 566.9500 639.8000 567.0500 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 542.9500 639.8000 543.0500 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 518.9500 639.8000 519.0500 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 494.9500 639.8000 495.0500 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 470.9500 639.8000 471.0500 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 446.9500 639.8000 447.0500 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 422.9500 639.8000 423.0500 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 398.9500 639.8000 399.0500 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 374.9500 639.8000 375.0500 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 350.9500 639.8000 351.0500 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 326.9500 639.8000 327.0500 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 302.9500 639.8000 303.0500 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 278.9500 639.8000 279.0500 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 254.9500 639.8000 255.0500 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 230.9500 639.8000 231.0500 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 206.9500 639.8000 207.0500 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 182.9500 639.8000 183.0500 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 158.9500 639.8000 159.0500 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 134.9500 639.8000 135.0500 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 110.9500 639.8000 111.0500 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 86.9500 639.8000 87.0500 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 62.9500 639.8000 63.0500 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 38.9500 639.8000 39.0500 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 639.2800 14.9500 639.8000 15.0500 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 249.3500 0.5200 249.4500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 245.5500 0.5200 245.6500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 241.7500 0.5200 241.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 237.9500 0.5200 238.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 234.1500 0.5200 234.2500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 230.3500 0.5200 230.4500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 226.5500 0.5200 226.6500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 222.7500 0.5200 222.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 218.9500 0.5200 219.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 215.1500 0.5200 215.2500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 211.3500 0.5200 211.4500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 207.5500 0.5200 207.6500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 203.7500 0.5200 203.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 199.9500 0.5200 200.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 196.1500 0.5200 196.2500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 192.3500 0.5200 192.4500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 188.5500 0.5200 188.6500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 184.7500 0.5200 184.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 180.9500 0.5200 181.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 177.1500 0.5200 177.2500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 173.3500 0.5200 173.4500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 169.5500 0.5200 169.6500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 165.7500 0.5200 165.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 161.9500 0.5200 162.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 158.1500 0.5200 158.2500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 154.3500 0.5200 154.4500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 150.5500 0.5200 150.6500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 146.7500 0.5200 146.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 142.9500 0.5200 143.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 139.1500 0.5200 139.2500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 135.3500 0.5200 135.4500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 131.5500 0.5200 131.6500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 127.7500 0.5200 127.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 123.9500 0.5200 124.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 120.1500 0.5200 120.2500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 116.3500 0.5200 116.4500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 112.5500 0.5200 112.6500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 108.7500 0.5200 108.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 104.9500 0.5200 105.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 101.1500 0.5200 101.2500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 97.3500 0.5200 97.4500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 93.5500 0.5200 93.6500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 89.7500 0.5200 89.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 85.9500 0.5200 86.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 82.1500 0.5200 82.2500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 78.3500 0.5200 78.4500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 74.5500 0.5200 74.6500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 70.7500 0.5200 70.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 66.9500 0.5200 67.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 63.1500 0.5200 63.2500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 59.3500 0.5200 59.4500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 55.5500 0.5200 55.6500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 51.7500 0.5200 51.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 47.9500 0.5200 48.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 44.1500 0.5200 44.2500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 40.3500 0.5200 40.4500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 36.5500 0.5200 36.6500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 32.7500 0.5200 32.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 28.9500 0.5200 29.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 25.1500 0.5200 25.2500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 21.3500 0.5200 21.4500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 17.5500 0.5200 17.6500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 13.7500 0.5200 13.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 9.9500 0.5200 10.0500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 571.4500 0.0000 571.5500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 564.4500 0.0000 564.5500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 557.4500 0.0000 557.5500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 550.4500 0.0000 550.5500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 543.4500 0.0000 543.5500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 536.4500 0.0000 536.5500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 529.4500 0.0000 529.5500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 522.4500 0.0000 522.5500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 515.4500 0.0000 515.5500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 508.4500 0.0000 508.5500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 501.4500 0.0000 501.5500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 494.4500 0.0000 494.5500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 487.4500 0.0000 487.5500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 480.4500 0.0000 480.5500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 473.4500 0.0000 473.5500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 466.4500 0.0000 466.5500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 459.4500 0.0000 459.5500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 452.4500 0.0000 452.5500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 445.4500 0.0000 445.5500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 438.4500 0.0000 438.5500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 431.4500 0.0000 431.5500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 424.4500 0.0000 424.5500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 417.4500 0.0000 417.5500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 410.4500 0.0000 410.5500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 403.4500 0.0000 403.5500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 396.4500 0.0000 396.5500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 389.4500 0.0000 389.5500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 382.4500 0.0000 382.5500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 375.4500 0.0000 375.5500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 368.4500 0.0000 368.5500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 361.4500 0.0000 361.5500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 354.4500 0.0000 354.5500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 347.4500 0.0000 347.5500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 340.4500 0.0000 340.5500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 333.4500 0.0000 333.5500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 326.4500 0.0000 326.5500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 319.4500 0.0000 319.5500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 312.4500 0.0000 312.5500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 305.4500 0.0000 305.5500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 298.4500 0.0000 298.5500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 291.4500 0.0000 291.5500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 284.4500 0.0000 284.5500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 277.4500 0.0000 277.5500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 270.4500 0.0000 270.5500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 263.4500 0.0000 263.5500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 256.4500 0.0000 256.5500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 249.4500 0.0000 249.5500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 242.4500 0.0000 242.5500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 235.4500 0.0000 235.5500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 228.4500 0.0000 228.5500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 221.4500 0.0000 221.5500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 214.4500 0.0000 214.5500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 207.4500 0.0000 207.5500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 200.4500 0.0000 200.5500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 193.4500 0.0000 193.5500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 186.4500 0.0000 186.5500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 179.4500 0.0000 179.5500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 172.4500 0.0000 172.5500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 165.4500 0.0000 165.5500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 158.4500 0.0000 158.5500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 151.4500 0.0000 151.5500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 144.4500 0.0000 144.5500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 137.4500 0.0000 137.5500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 130.4500 0.0000 130.5500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 123.4500 0.0000 123.5500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 116.4500 0.0000 116.5500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 109.4500 0.0000 109.5500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 102.4500 0.0000 102.5500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 95.4500 0.0000 95.5500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 88.4500 0.0000 88.5500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 81.4500 0.0000 81.5500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 74.4500 0.0000 74.5500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 67.4500 0.0000 67.5500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 60.4500 0.0000 60.5500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 53.4500 0.0000 53.5500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 46.4500 0.0000 46.5500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 39.4500 0.0000 39.5500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 32.4500 0.0000 32.5500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 25.4500 0.0000 25.5500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 18.4500 0.0000 18.5500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 568.0500 0.0000 568.1500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 561.0500 0.0000 561.1500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.0500 0.0000 554.1500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 547.0500 0.0000 547.1500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 540.0500 0.0000 540.1500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 533.0500 0.0000 533.1500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 526.0500 0.0000 526.1500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 519.0500 0.0000 519.1500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 512.0500 0.0000 512.1500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 505.0500 0.0000 505.1500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.0500 0.0000 498.1500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 491.0500 0.0000 491.1500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 484.0500 0.0000 484.1500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 477.0500 0.0000 477.1500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.0500 0.0000 470.1500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 463.0500 0.0000 463.1500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 456.0500 0.0000 456.1500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 449.0500 0.0000 449.1500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 442.0500 0.0000 442.1500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 435.0500 0.0000 435.1500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 428.0500 0.0000 428.1500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 421.0500 0.0000 421.1500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 414.0500 0.0000 414.1500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 407.0500 0.0000 407.1500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 400.0500 0.0000 400.1500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 393.0500 0.0000 393.1500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 386.0500 0.0000 386.1500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 379.0500 0.0000 379.1500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 372.0500 0.0000 372.1500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 365.0500 0.0000 365.1500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 358.0500 0.0000 358.1500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 351.0500 0.0000 351.1500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 344.0500 0.0000 344.1500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 337.0500 0.0000 337.1500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 330.0500 0.0000 330.1500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 323.0500 0.0000 323.1500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 316.0500 0.0000 316.1500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 309.0500 0.0000 309.1500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 302.0500 0.0000 302.1500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 295.0500 0.0000 295.1500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 288.0500 0.0000 288.1500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 281.0500 0.0000 281.1500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 274.0500 0.0000 274.1500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 267.0500 0.0000 267.1500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 260.0500 0.0000 260.1500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 253.0500 0.0000 253.1500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 246.0500 0.0000 246.1500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 239.0500 0.0000 239.1500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 232.0500 0.0000 232.1500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 225.0500 0.0000 225.1500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 218.0500 0.0000 218.1500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 211.0500 0.0000 211.1500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 204.0500 0.0000 204.1500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 197.0500 0.0000 197.1500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 190.0500 0.0000 190.1500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 183.0500 0.0000 183.1500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 176.0500 0.0000 176.1500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 169.0500 0.0000 169.1500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 162.0500 0.0000 162.1500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 155.0500 0.0000 155.1500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 148.0500 0.0000 148.1500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 141.0500 0.0000 141.1500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 134.0500 0.0000 134.1500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 127.0500 0.0000 127.1500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 120.0500 0.0000 120.1500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 113.0500 0.0000 113.1500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 106.0500 0.0000 106.1500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 99.0500 0.0000 99.1500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 92.0500 0.0000 92.1500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 85.0500 0.0000 85.1500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 78.0500 0.0000 78.1500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 71.0500 0.0000 71.1500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 64.0500 0.0000 64.1500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.0500 0.0000 57.1500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 50.0500 0.0000 50.1500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 43.0500 0.0000 43.1500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 36.0500 0.0000 36.1500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 29.0500 0.0000 29.1500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 22.0500 0.0000 22.1500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 15.0500 0.0000 15.1500 0.5200 ;
    END
  END out[0]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 321.5500 0.5200 321.6500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 317.7500 0.5200 317.8500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 313.9500 0.5200 314.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 310.1500 0.5200 310.2500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 306.3500 0.5200 306.4500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 302.5500 0.5200 302.6500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 298.7500 0.5200 298.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 294.9500 0.5200 295.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 291.1500 0.5200 291.2500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 287.3500 0.5200 287.4500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 283.5500 0.5200 283.6500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 279.7500 0.5200 279.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 275.9500 0.5200 276.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 272.1500 0.5200 272.2500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 268.3500 0.5200 268.4500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 264.5500 0.5200 264.6500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 260.7500 0.5200 260.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 256.9500 0.5200 257.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 253.1500 0.5200 253.2500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 329.1500 0.5200 329.2500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 639.8000 639.2000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 639.8000 639.2000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 639.8000 639.2000 ;
    LAYER M4 ;
      RECT 0.0000 0.6200 639.8000 639.2000 ;
      RECT 568.2500 0.0000 639.8000 0.6200 ;
      RECT 561.2500 0.0000 567.9500 0.6200 ;
      RECT 554.2500 0.0000 560.9500 0.6200 ;
      RECT 547.2500 0.0000 553.9500 0.6200 ;
      RECT 540.2500 0.0000 546.9500 0.6200 ;
      RECT 533.2500 0.0000 539.9500 0.6200 ;
      RECT 526.2500 0.0000 532.9500 0.6200 ;
      RECT 519.2500 0.0000 525.9500 0.6200 ;
      RECT 512.2500 0.0000 518.9500 0.6200 ;
      RECT 505.2500 0.0000 511.9500 0.6200 ;
      RECT 498.2500 0.0000 504.9500 0.6200 ;
      RECT 491.2500 0.0000 497.9500 0.6200 ;
      RECT 484.2500 0.0000 490.9500 0.6200 ;
      RECT 477.2500 0.0000 483.9500 0.6200 ;
      RECT 470.2500 0.0000 476.9500 0.6200 ;
      RECT 463.2500 0.0000 469.9500 0.6200 ;
      RECT 456.2500 0.0000 462.9500 0.6200 ;
      RECT 449.2500 0.0000 455.9500 0.6200 ;
      RECT 442.2500 0.0000 448.9500 0.6200 ;
      RECT 435.2500 0.0000 441.9500 0.6200 ;
      RECT 428.2500 0.0000 434.9500 0.6200 ;
      RECT 421.2500 0.0000 427.9500 0.6200 ;
      RECT 414.2500 0.0000 420.9500 0.6200 ;
      RECT 407.2500 0.0000 413.9500 0.6200 ;
      RECT 400.2500 0.0000 406.9500 0.6200 ;
      RECT 393.2500 0.0000 399.9500 0.6200 ;
      RECT 386.2500 0.0000 392.9500 0.6200 ;
      RECT 379.2500 0.0000 385.9500 0.6200 ;
      RECT 372.2500 0.0000 378.9500 0.6200 ;
      RECT 365.2500 0.0000 371.9500 0.6200 ;
      RECT 358.2500 0.0000 364.9500 0.6200 ;
      RECT 351.2500 0.0000 357.9500 0.6200 ;
      RECT 344.2500 0.0000 350.9500 0.6200 ;
      RECT 337.2500 0.0000 343.9500 0.6200 ;
      RECT 330.2500 0.0000 336.9500 0.6200 ;
      RECT 323.2500 0.0000 329.9500 0.6200 ;
      RECT 316.2500 0.0000 322.9500 0.6200 ;
      RECT 309.2500 0.0000 315.9500 0.6200 ;
      RECT 302.2500 0.0000 308.9500 0.6200 ;
      RECT 295.2500 0.0000 301.9500 0.6200 ;
      RECT 288.2500 0.0000 294.9500 0.6200 ;
      RECT 281.2500 0.0000 287.9500 0.6200 ;
      RECT 274.2500 0.0000 280.9500 0.6200 ;
      RECT 267.2500 0.0000 273.9500 0.6200 ;
      RECT 260.2500 0.0000 266.9500 0.6200 ;
      RECT 253.2500 0.0000 259.9500 0.6200 ;
      RECT 246.2500 0.0000 252.9500 0.6200 ;
      RECT 239.2500 0.0000 245.9500 0.6200 ;
      RECT 232.2500 0.0000 238.9500 0.6200 ;
      RECT 225.2500 0.0000 231.9500 0.6200 ;
      RECT 218.2500 0.0000 224.9500 0.6200 ;
      RECT 211.2500 0.0000 217.9500 0.6200 ;
      RECT 204.2500 0.0000 210.9500 0.6200 ;
      RECT 197.2500 0.0000 203.9500 0.6200 ;
      RECT 190.2500 0.0000 196.9500 0.6200 ;
      RECT 183.2500 0.0000 189.9500 0.6200 ;
      RECT 176.2500 0.0000 182.9500 0.6200 ;
      RECT 169.2500 0.0000 175.9500 0.6200 ;
      RECT 162.2500 0.0000 168.9500 0.6200 ;
      RECT 155.2500 0.0000 161.9500 0.6200 ;
      RECT 148.2500 0.0000 154.9500 0.6200 ;
      RECT 141.2500 0.0000 147.9500 0.6200 ;
      RECT 134.2500 0.0000 140.9500 0.6200 ;
      RECT 127.2500 0.0000 133.9500 0.6200 ;
      RECT 120.2500 0.0000 126.9500 0.6200 ;
      RECT 113.2500 0.0000 119.9500 0.6200 ;
      RECT 106.2500 0.0000 112.9500 0.6200 ;
      RECT 99.2500 0.0000 105.9500 0.6200 ;
      RECT 92.2500 0.0000 98.9500 0.6200 ;
      RECT 85.2500 0.0000 91.9500 0.6200 ;
      RECT 78.2500 0.0000 84.9500 0.6200 ;
      RECT 71.2500 0.0000 77.9500 0.6200 ;
      RECT 64.2500 0.0000 70.9500 0.6200 ;
      RECT 57.2500 0.0000 63.9500 0.6200 ;
      RECT 50.2500 0.0000 56.9500 0.6200 ;
      RECT 43.2500 0.0000 49.9500 0.6200 ;
      RECT 36.2500 0.0000 42.9500 0.6200 ;
      RECT 29.2500 0.0000 35.9500 0.6200 ;
      RECT 22.2500 0.0000 28.9500 0.6200 ;
      RECT 15.2500 0.0000 21.9500 0.6200 ;
      RECT 0.0000 0.0000 14.9500 0.6200 ;
    LAYER M5 ;
      RECT 0.0000 567.1500 639.8000 639.2000 ;
      RECT 0.0000 566.8500 639.1800 567.1500 ;
      RECT 0.0000 543.1500 639.8000 566.8500 ;
      RECT 0.0000 542.8500 639.1800 543.1500 ;
      RECT 0.0000 519.1500 639.8000 542.8500 ;
      RECT 0.0000 518.8500 639.1800 519.1500 ;
      RECT 0.0000 495.1500 639.8000 518.8500 ;
      RECT 0.0000 494.8500 639.1800 495.1500 ;
      RECT 0.0000 471.1500 639.8000 494.8500 ;
      RECT 0.0000 470.8500 639.1800 471.1500 ;
      RECT 0.0000 447.1500 639.8000 470.8500 ;
      RECT 0.0000 446.8500 639.1800 447.1500 ;
      RECT 0.0000 423.1500 639.8000 446.8500 ;
      RECT 0.0000 422.8500 639.1800 423.1500 ;
      RECT 0.0000 399.1500 639.8000 422.8500 ;
      RECT 0.0000 398.8500 639.1800 399.1500 ;
      RECT 0.0000 375.1500 639.8000 398.8500 ;
      RECT 0.0000 374.8500 639.1800 375.1500 ;
      RECT 0.0000 351.1500 639.8000 374.8500 ;
      RECT 0.0000 350.8500 639.1800 351.1500 ;
      RECT 0.0000 329.3500 639.8000 350.8500 ;
      RECT 0.6200 329.0500 639.8000 329.3500 ;
      RECT 0.0000 327.1500 639.8000 329.0500 ;
      RECT 0.0000 326.8500 639.1800 327.1500 ;
      RECT 0.0000 325.5500 639.8000 326.8500 ;
      RECT 0.6200 325.2500 639.8000 325.5500 ;
      RECT 0.0000 321.7500 639.8000 325.2500 ;
      RECT 0.6200 321.4500 639.8000 321.7500 ;
      RECT 0.0000 317.9500 639.8000 321.4500 ;
      RECT 0.6200 317.6500 639.8000 317.9500 ;
      RECT 0.0000 314.1500 639.8000 317.6500 ;
      RECT 0.6200 313.8500 639.8000 314.1500 ;
      RECT 0.0000 310.3500 639.8000 313.8500 ;
      RECT 0.6200 310.0500 639.8000 310.3500 ;
      RECT 0.0000 306.5500 639.8000 310.0500 ;
      RECT 0.6200 306.2500 639.8000 306.5500 ;
      RECT 0.0000 303.1500 639.8000 306.2500 ;
      RECT 0.0000 302.8500 639.1800 303.1500 ;
      RECT 0.0000 302.7500 639.8000 302.8500 ;
      RECT 0.6200 302.4500 639.8000 302.7500 ;
      RECT 0.0000 298.9500 639.8000 302.4500 ;
      RECT 0.6200 298.6500 639.8000 298.9500 ;
      RECT 0.0000 295.1500 639.8000 298.6500 ;
      RECT 0.6200 294.8500 639.8000 295.1500 ;
      RECT 0.0000 291.3500 639.8000 294.8500 ;
      RECT 0.6200 291.0500 639.8000 291.3500 ;
      RECT 0.0000 287.5500 639.8000 291.0500 ;
      RECT 0.6200 287.2500 639.8000 287.5500 ;
      RECT 0.0000 283.7500 639.8000 287.2500 ;
      RECT 0.6200 283.4500 639.8000 283.7500 ;
      RECT 0.0000 279.9500 639.8000 283.4500 ;
      RECT 0.6200 279.6500 639.8000 279.9500 ;
      RECT 0.0000 279.1500 639.8000 279.6500 ;
      RECT 0.0000 278.8500 639.1800 279.1500 ;
      RECT 0.0000 276.1500 639.8000 278.8500 ;
      RECT 0.6200 275.8500 639.8000 276.1500 ;
      RECT 0.0000 272.3500 639.8000 275.8500 ;
      RECT 0.6200 272.0500 639.8000 272.3500 ;
      RECT 0.0000 268.5500 639.8000 272.0500 ;
      RECT 0.6200 268.2500 639.8000 268.5500 ;
      RECT 0.0000 264.7500 639.8000 268.2500 ;
      RECT 0.6200 264.4500 639.8000 264.7500 ;
      RECT 0.0000 260.9500 639.8000 264.4500 ;
      RECT 0.6200 260.6500 639.8000 260.9500 ;
      RECT 0.0000 257.1500 639.8000 260.6500 ;
      RECT 0.6200 256.8500 639.8000 257.1500 ;
      RECT 0.0000 255.1500 639.8000 256.8500 ;
      RECT 0.0000 254.8500 639.1800 255.1500 ;
      RECT 0.0000 253.3500 639.8000 254.8500 ;
      RECT 0.6200 253.0500 639.8000 253.3500 ;
      RECT 0.0000 249.5500 639.8000 253.0500 ;
      RECT 0.6200 249.2500 639.8000 249.5500 ;
      RECT 0.0000 245.7500 639.8000 249.2500 ;
      RECT 0.6200 245.4500 639.8000 245.7500 ;
      RECT 0.0000 241.9500 639.8000 245.4500 ;
      RECT 0.6200 241.6500 639.8000 241.9500 ;
      RECT 0.0000 238.1500 639.8000 241.6500 ;
      RECT 0.6200 237.8500 639.8000 238.1500 ;
      RECT 0.0000 234.3500 639.8000 237.8500 ;
      RECT 0.6200 234.0500 639.8000 234.3500 ;
      RECT 0.0000 231.1500 639.8000 234.0500 ;
      RECT 0.0000 230.8500 639.1800 231.1500 ;
      RECT 0.0000 230.5500 639.8000 230.8500 ;
      RECT 0.6200 230.2500 639.8000 230.5500 ;
      RECT 0.0000 226.7500 639.8000 230.2500 ;
      RECT 0.6200 226.4500 639.8000 226.7500 ;
      RECT 0.0000 222.9500 639.8000 226.4500 ;
      RECT 0.6200 222.6500 639.8000 222.9500 ;
      RECT 0.0000 219.1500 639.8000 222.6500 ;
      RECT 0.6200 218.8500 639.8000 219.1500 ;
      RECT 0.0000 215.3500 639.8000 218.8500 ;
      RECT 0.6200 215.0500 639.8000 215.3500 ;
      RECT 0.0000 211.5500 639.8000 215.0500 ;
      RECT 0.6200 211.2500 639.8000 211.5500 ;
      RECT 0.0000 207.7500 639.8000 211.2500 ;
      RECT 0.6200 207.4500 639.8000 207.7500 ;
      RECT 0.0000 207.1500 639.8000 207.4500 ;
      RECT 0.0000 206.8500 639.1800 207.1500 ;
      RECT 0.0000 203.9500 639.8000 206.8500 ;
      RECT 0.6200 203.6500 639.8000 203.9500 ;
      RECT 0.0000 200.1500 639.8000 203.6500 ;
      RECT 0.6200 199.8500 639.8000 200.1500 ;
      RECT 0.0000 196.3500 639.8000 199.8500 ;
      RECT 0.6200 196.0500 639.8000 196.3500 ;
      RECT 0.0000 192.5500 639.8000 196.0500 ;
      RECT 0.6200 192.2500 639.8000 192.5500 ;
      RECT 0.0000 188.7500 639.8000 192.2500 ;
      RECT 0.6200 188.4500 639.8000 188.7500 ;
      RECT 0.0000 184.9500 639.8000 188.4500 ;
      RECT 0.6200 184.6500 639.8000 184.9500 ;
      RECT 0.0000 183.1500 639.8000 184.6500 ;
      RECT 0.0000 182.8500 639.1800 183.1500 ;
      RECT 0.0000 181.1500 639.8000 182.8500 ;
      RECT 0.6200 180.8500 639.8000 181.1500 ;
      RECT 0.0000 177.3500 639.8000 180.8500 ;
      RECT 0.6200 177.0500 639.8000 177.3500 ;
      RECT 0.0000 173.5500 639.8000 177.0500 ;
      RECT 0.6200 173.2500 639.8000 173.5500 ;
      RECT 0.0000 169.7500 639.8000 173.2500 ;
      RECT 0.6200 169.4500 639.8000 169.7500 ;
      RECT 0.0000 165.9500 639.8000 169.4500 ;
      RECT 0.6200 165.6500 639.8000 165.9500 ;
      RECT 0.0000 162.1500 639.8000 165.6500 ;
      RECT 0.6200 161.8500 639.8000 162.1500 ;
      RECT 0.0000 159.1500 639.8000 161.8500 ;
      RECT 0.0000 158.8500 639.1800 159.1500 ;
      RECT 0.0000 158.3500 639.8000 158.8500 ;
      RECT 0.6200 158.0500 639.8000 158.3500 ;
      RECT 0.0000 154.5500 639.8000 158.0500 ;
      RECT 0.6200 154.2500 639.8000 154.5500 ;
      RECT 0.0000 150.7500 639.8000 154.2500 ;
      RECT 0.6200 150.4500 639.8000 150.7500 ;
      RECT 0.0000 146.9500 639.8000 150.4500 ;
      RECT 0.6200 146.6500 639.8000 146.9500 ;
      RECT 0.0000 143.1500 639.8000 146.6500 ;
      RECT 0.6200 142.8500 639.8000 143.1500 ;
      RECT 0.0000 139.3500 639.8000 142.8500 ;
      RECT 0.6200 139.0500 639.8000 139.3500 ;
      RECT 0.0000 135.5500 639.8000 139.0500 ;
      RECT 0.6200 135.2500 639.8000 135.5500 ;
      RECT 0.0000 135.1500 639.8000 135.2500 ;
      RECT 0.0000 134.8500 639.1800 135.1500 ;
      RECT 0.0000 131.7500 639.8000 134.8500 ;
      RECT 0.6200 131.4500 639.8000 131.7500 ;
      RECT 0.0000 127.9500 639.8000 131.4500 ;
      RECT 0.6200 127.6500 639.8000 127.9500 ;
      RECT 0.0000 124.1500 639.8000 127.6500 ;
      RECT 0.6200 123.8500 639.8000 124.1500 ;
      RECT 0.0000 120.3500 639.8000 123.8500 ;
      RECT 0.6200 120.0500 639.8000 120.3500 ;
      RECT 0.0000 116.5500 639.8000 120.0500 ;
      RECT 0.6200 116.2500 639.8000 116.5500 ;
      RECT 0.0000 112.7500 639.8000 116.2500 ;
      RECT 0.6200 112.4500 639.8000 112.7500 ;
      RECT 0.0000 111.1500 639.8000 112.4500 ;
      RECT 0.0000 110.8500 639.1800 111.1500 ;
      RECT 0.0000 108.9500 639.8000 110.8500 ;
      RECT 0.6200 108.6500 639.8000 108.9500 ;
      RECT 0.0000 105.1500 639.8000 108.6500 ;
      RECT 0.6200 104.8500 639.8000 105.1500 ;
      RECT 0.0000 101.3500 639.8000 104.8500 ;
      RECT 0.6200 101.0500 639.8000 101.3500 ;
      RECT 0.0000 97.5500 639.8000 101.0500 ;
      RECT 0.6200 97.2500 639.8000 97.5500 ;
      RECT 0.0000 93.7500 639.8000 97.2500 ;
      RECT 0.6200 93.4500 639.8000 93.7500 ;
      RECT 0.0000 89.9500 639.8000 93.4500 ;
      RECT 0.6200 89.6500 639.8000 89.9500 ;
      RECT 0.0000 87.1500 639.8000 89.6500 ;
      RECT 0.0000 86.8500 639.1800 87.1500 ;
      RECT 0.0000 86.1500 639.8000 86.8500 ;
      RECT 0.6200 85.8500 639.8000 86.1500 ;
      RECT 0.0000 82.3500 639.8000 85.8500 ;
      RECT 0.6200 82.0500 639.8000 82.3500 ;
      RECT 0.0000 78.5500 639.8000 82.0500 ;
      RECT 0.6200 78.2500 639.8000 78.5500 ;
      RECT 0.0000 74.7500 639.8000 78.2500 ;
      RECT 0.6200 74.4500 639.8000 74.7500 ;
      RECT 0.0000 70.9500 639.8000 74.4500 ;
      RECT 0.6200 70.6500 639.8000 70.9500 ;
      RECT 0.0000 67.1500 639.8000 70.6500 ;
      RECT 0.6200 66.8500 639.8000 67.1500 ;
      RECT 0.0000 63.3500 639.8000 66.8500 ;
      RECT 0.6200 63.1500 639.8000 63.3500 ;
      RECT 0.6200 63.0500 639.1800 63.1500 ;
      RECT 0.0000 62.8500 639.1800 63.0500 ;
      RECT 0.0000 59.5500 639.8000 62.8500 ;
      RECT 0.6200 59.2500 639.8000 59.5500 ;
      RECT 0.0000 55.7500 639.8000 59.2500 ;
      RECT 0.6200 55.4500 639.8000 55.7500 ;
      RECT 0.0000 51.9500 639.8000 55.4500 ;
      RECT 0.6200 51.6500 639.8000 51.9500 ;
      RECT 0.0000 48.1500 639.8000 51.6500 ;
      RECT 0.6200 47.8500 639.8000 48.1500 ;
      RECT 0.0000 44.3500 639.8000 47.8500 ;
      RECT 0.6200 44.0500 639.8000 44.3500 ;
      RECT 0.0000 40.5500 639.8000 44.0500 ;
      RECT 0.6200 40.2500 639.8000 40.5500 ;
      RECT 0.0000 39.1500 639.8000 40.2500 ;
      RECT 0.0000 38.8500 639.1800 39.1500 ;
      RECT 0.0000 36.7500 639.8000 38.8500 ;
      RECT 0.6200 36.4500 639.8000 36.7500 ;
      RECT 0.0000 32.9500 639.8000 36.4500 ;
      RECT 0.6200 32.6500 639.8000 32.9500 ;
      RECT 0.0000 29.1500 639.8000 32.6500 ;
      RECT 0.6200 28.8500 639.8000 29.1500 ;
      RECT 0.0000 25.3500 639.8000 28.8500 ;
      RECT 0.6200 25.0500 639.8000 25.3500 ;
      RECT 0.0000 21.5500 639.8000 25.0500 ;
      RECT 0.6200 21.2500 639.8000 21.5500 ;
      RECT 0.0000 17.7500 639.8000 21.2500 ;
      RECT 0.6200 17.4500 639.8000 17.7500 ;
      RECT 0.0000 15.1500 639.8000 17.4500 ;
      RECT 0.0000 14.8500 639.1800 15.1500 ;
      RECT 0.0000 13.9500 639.8000 14.8500 ;
      RECT 0.6200 13.6500 639.8000 13.9500 ;
      RECT 0.0000 10.1500 639.8000 13.6500 ;
      RECT 0.6200 9.8500 639.8000 10.1500 ;
      RECT 0.0000 0.0000 639.8000 9.8500 ;
    LAYER M6 ;
      RECT 0.0000 0.6200 639.8000 639.2000 ;
      RECT 571.6500 0.0000 639.8000 0.6200 ;
      RECT 564.6500 0.0000 571.3500 0.6200 ;
      RECT 557.6500 0.0000 564.3500 0.6200 ;
      RECT 550.6500 0.0000 557.3500 0.6200 ;
      RECT 543.6500 0.0000 550.3500 0.6200 ;
      RECT 536.6500 0.0000 543.3500 0.6200 ;
      RECT 529.6500 0.0000 536.3500 0.6200 ;
      RECT 522.6500 0.0000 529.3500 0.6200 ;
      RECT 515.6500 0.0000 522.3500 0.6200 ;
      RECT 508.6500 0.0000 515.3500 0.6200 ;
      RECT 501.6500 0.0000 508.3500 0.6200 ;
      RECT 494.6500 0.0000 501.3500 0.6200 ;
      RECT 487.6500 0.0000 494.3500 0.6200 ;
      RECT 480.6500 0.0000 487.3500 0.6200 ;
      RECT 473.6500 0.0000 480.3500 0.6200 ;
      RECT 466.6500 0.0000 473.3500 0.6200 ;
      RECT 459.6500 0.0000 466.3500 0.6200 ;
      RECT 452.6500 0.0000 459.3500 0.6200 ;
      RECT 445.6500 0.0000 452.3500 0.6200 ;
      RECT 438.6500 0.0000 445.3500 0.6200 ;
      RECT 431.6500 0.0000 438.3500 0.6200 ;
      RECT 424.6500 0.0000 431.3500 0.6200 ;
      RECT 417.6500 0.0000 424.3500 0.6200 ;
      RECT 410.6500 0.0000 417.3500 0.6200 ;
      RECT 403.6500 0.0000 410.3500 0.6200 ;
      RECT 396.6500 0.0000 403.3500 0.6200 ;
      RECT 389.6500 0.0000 396.3500 0.6200 ;
      RECT 382.6500 0.0000 389.3500 0.6200 ;
      RECT 375.6500 0.0000 382.3500 0.6200 ;
      RECT 368.6500 0.0000 375.3500 0.6200 ;
      RECT 361.6500 0.0000 368.3500 0.6200 ;
      RECT 354.6500 0.0000 361.3500 0.6200 ;
      RECT 347.6500 0.0000 354.3500 0.6200 ;
      RECT 340.6500 0.0000 347.3500 0.6200 ;
      RECT 333.6500 0.0000 340.3500 0.6200 ;
      RECT 326.6500 0.0000 333.3500 0.6200 ;
      RECT 319.6500 0.0000 326.3500 0.6200 ;
      RECT 312.6500 0.0000 319.3500 0.6200 ;
      RECT 305.6500 0.0000 312.3500 0.6200 ;
      RECT 298.6500 0.0000 305.3500 0.6200 ;
      RECT 291.6500 0.0000 298.3500 0.6200 ;
      RECT 284.6500 0.0000 291.3500 0.6200 ;
      RECT 277.6500 0.0000 284.3500 0.6200 ;
      RECT 270.6500 0.0000 277.3500 0.6200 ;
      RECT 263.6500 0.0000 270.3500 0.6200 ;
      RECT 256.6500 0.0000 263.3500 0.6200 ;
      RECT 249.6500 0.0000 256.3500 0.6200 ;
      RECT 242.6500 0.0000 249.3500 0.6200 ;
      RECT 235.6500 0.0000 242.3500 0.6200 ;
      RECT 228.6500 0.0000 235.3500 0.6200 ;
      RECT 221.6500 0.0000 228.3500 0.6200 ;
      RECT 214.6500 0.0000 221.3500 0.6200 ;
      RECT 207.6500 0.0000 214.3500 0.6200 ;
      RECT 200.6500 0.0000 207.3500 0.6200 ;
      RECT 193.6500 0.0000 200.3500 0.6200 ;
      RECT 186.6500 0.0000 193.3500 0.6200 ;
      RECT 179.6500 0.0000 186.3500 0.6200 ;
      RECT 172.6500 0.0000 179.3500 0.6200 ;
      RECT 165.6500 0.0000 172.3500 0.6200 ;
      RECT 158.6500 0.0000 165.3500 0.6200 ;
      RECT 151.6500 0.0000 158.3500 0.6200 ;
      RECT 144.6500 0.0000 151.3500 0.6200 ;
      RECT 137.6500 0.0000 144.3500 0.6200 ;
      RECT 130.6500 0.0000 137.3500 0.6200 ;
      RECT 123.6500 0.0000 130.3500 0.6200 ;
      RECT 116.6500 0.0000 123.3500 0.6200 ;
      RECT 109.6500 0.0000 116.3500 0.6200 ;
      RECT 102.6500 0.0000 109.3500 0.6200 ;
      RECT 95.6500 0.0000 102.3500 0.6200 ;
      RECT 88.6500 0.0000 95.3500 0.6200 ;
      RECT 81.6500 0.0000 88.3500 0.6200 ;
      RECT 74.6500 0.0000 81.3500 0.6200 ;
      RECT 67.6500 0.0000 74.3500 0.6200 ;
      RECT 60.6500 0.0000 67.3500 0.6200 ;
      RECT 53.6500 0.0000 60.3500 0.6200 ;
      RECT 46.6500 0.0000 53.3500 0.6200 ;
      RECT 39.6500 0.0000 46.3500 0.6200 ;
      RECT 32.6500 0.0000 39.3500 0.6200 ;
      RECT 25.6500 0.0000 32.3500 0.6200 ;
      RECT 18.6500 0.0000 25.3500 0.6200 ;
      RECT 0.0000 0.0000 18.3500 0.6200 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 639.8000 639.2000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 639.8000 639.2000 ;
  END
END core

END LIBRARY
