##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar  8 16:42:16 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w8
  CLASS BLOCK ;
  SIZE 163.8000 BY 160.6000 ;
  FOREIGN sram_w8 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 68.3500 0.6000 68.4500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.0500 0.0000 145.1500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.0500 0.0000 144.1500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.0500 0.0000 143.1500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.0500 0.0000 142.1500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.0500 0.0000 141.1500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.0500 0.0000 140.1500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.0500 0.0000 139.1500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.0500 0.0000 138.1500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 0.0000 137.1500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.0500 0.0000 136.1500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.0500 0.0000 135.1500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 0.0000 134.1500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 0.0000 133.1500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.0500 0.0000 132.1500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.0500 0.0000 131.1500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.0500 0.0000 130.1500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.0500 0.0000 129.1500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.0500 0.0000 128.1500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.0500 0.0000 127.1500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 0.0000 126.1500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.0500 0.0000 125.1500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0500 0.0000 124.1500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.0500 0.0000 123.1500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.0500 0.0000 122.1500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 0.0000 121.1500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.0500 0.0000 120.1500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 0.0000 119.1500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.0500 0.0000 118.1500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.0500 0.0000 117.1500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.0500 0.0000 116.1500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.0500 0.0000 115.1500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.0500 0.0000 114.1500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.0500 0.0000 113.1500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.0500 0.0000 112.1500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 0.0000 111.1500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 0.0000 110.1500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 0.0000 109.1500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.0500 0.0000 108.1500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.0500 0.0000 107.1500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 0.0000 106.1500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.0500 0.0000 105.1500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.0500 0.0000 104.1500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.0500 0.0000 103.1500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 0.0000 102.1500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 0.0000 101.1500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.0500 0.0000 100.1500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.0500 0.0000 99.1500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 0.0000 98.1500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.0500 0.0000 97.1500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.0500 0.0000 96.1500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.0500 0.0000 95.1500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 0.0000 94.1500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.0500 0.0000 93.1500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.0500 0.0000 92.1500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.0500 0.0000 91.1500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.0500 0.0000 90.1500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.0500 0.0000 89.1500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.0500 0.0000 88.1500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.0500 0.0000 87.1500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.0500 0.0000 86.1500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 0.0000 85.1500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.0500 0.0000 84.1500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.0500 0.0000 83.1500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.0500 0.0000 82.1500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.0500 0.0000 81.1500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.0500 0.0000 80.1500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.0500 0.0000 79.1500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.0500 0.0000 78.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.0500 0.0000 77.1500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.0500 0.0000 76.1500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.0500 0.0000 75.1500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 0.0000 74.1500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.0500 0.0000 73.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.0500 0.0000 72.1500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.0500 0.0000 71.1500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.0500 0.0000 70.1500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.0500 0.0000 69.1500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.0500 0.0000 68.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.0500 0.0000 67.1500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.0500 0.0000 66.1500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.0500 0.0000 65.1500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.0500 0.0000 64.1500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.0500 0.0000 63.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.0500 0.0000 62.1500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.0500 0.0000 61.1500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.0500 0.0000 60.1500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.0500 0.0000 59.1500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.0500 0.0000 58.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.0500 0.0000 57.1500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.0500 0.0000 56.1500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0500 0.0000 55.1500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.0500 0.0000 54.1500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.0500 0.0000 53.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.0500 0.0000 52.1500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.0500 0.0000 51.1500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.0500 0.0000 50.1500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.0500 0.0000 49.1500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.0500 0.0000 48.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.0500 0.0000 47.1500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0500 0.0000 46.1500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.0500 0.0000 45.1500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.0500 0.0000 44.1500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.0500 0.0000 43.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0500 0.0000 42.1500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.0500 0.0000 41.1500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.0500 0.0000 40.1500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.0500 0.0000 39.1500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0500 0.0000 38.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.0500 0.0000 37.1500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.0500 0.0000 36.1500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.0500 0.0000 35.1500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0500 0.0000 34.1500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0500 0.0000 33.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.0500 0.0000 32.1500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.0500 0.0000 31.1500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0500 0.0000 30.1500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0500 0.0000 29.1500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.0500 0.0000 28.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.0500 0.0000 27.1500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.0500 0.0000 26.1500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0500 0.0000 25.1500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.0500 0.0000 24.1500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.0500 0.0000 23.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.0500 0.0000 22.1500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0500 0.0000 21.1500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0500 0.0000 20.1500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.0500 0.0000 19.1500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 0.0000 18.1500 0.6000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.0500 160.0000 145.1500 160.6000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.0500 160.0000 144.1500 160.6000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.0500 160.0000 143.1500 160.6000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.0500 160.0000 142.1500 160.6000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.0500 160.0000 141.1500 160.6000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.0500 160.0000 140.1500 160.6000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.0500 160.0000 139.1500 160.6000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.0500 160.0000 138.1500 160.6000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.0500 160.0000 137.1500 160.6000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.0500 160.0000 136.1500 160.6000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.0500 160.0000 135.1500 160.6000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 160.0000 134.1500 160.6000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 160.0000 133.1500 160.6000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.0500 160.0000 132.1500 160.6000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.0500 160.0000 131.1500 160.6000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.0500 160.0000 130.1500 160.6000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.0500 160.0000 129.1500 160.6000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.0500 160.0000 128.1500 160.6000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.0500 160.0000 127.1500 160.6000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 160.0000 126.1500 160.6000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.0500 160.0000 125.1500 160.6000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0500 160.0000 124.1500 160.6000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.0500 160.0000 123.1500 160.6000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.0500 160.0000 122.1500 160.6000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 160.0000 121.1500 160.6000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.0500 160.0000 120.1500 160.6000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 160.0000 119.1500 160.6000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.0500 160.0000 118.1500 160.6000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.0500 160.0000 117.1500 160.6000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.0500 160.0000 116.1500 160.6000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.0500 160.0000 115.1500 160.6000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.0500 160.0000 114.1500 160.6000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.0500 160.0000 113.1500 160.6000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.0500 160.0000 112.1500 160.6000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 160.0000 111.1500 160.6000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 160.0000 110.1500 160.6000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 160.0000 109.1500 160.6000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.0500 160.0000 108.1500 160.6000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.0500 160.0000 107.1500 160.6000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 160.0000 106.1500 160.6000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.0500 160.0000 105.1500 160.6000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.0500 160.0000 104.1500 160.6000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.0500 160.0000 103.1500 160.6000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 160.0000 102.1500 160.6000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 160.0000 101.1500 160.6000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.0500 160.0000 100.1500 160.6000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.0500 160.0000 99.1500 160.6000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 160.0000 98.1500 160.6000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.0500 160.0000 97.1500 160.6000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.0500 160.0000 96.1500 160.6000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.0500 160.0000 95.1500 160.6000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 160.0000 94.1500 160.6000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.0500 160.0000 93.1500 160.6000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.0500 160.0000 92.1500 160.6000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.0500 160.0000 91.1500 160.6000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.0500 160.0000 90.1500 160.6000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.0500 160.0000 89.1500 160.6000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.0500 160.0000 88.1500 160.6000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.0500 160.0000 87.1500 160.6000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.0500 160.0000 86.1500 160.6000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.0500 160.0000 85.1500 160.6000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.0500 160.0000 84.1500 160.6000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.0500 160.0000 83.1500 160.6000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.0500 160.0000 82.1500 160.6000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.0500 160.0000 81.1500 160.6000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.0500 160.0000 80.1500 160.6000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.0500 160.0000 79.1500 160.6000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.0500 160.0000 78.1500 160.6000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.0500 160.0000 77.1500 160.6000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.0500 160.0000 76.1500 160.6000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.0500 160.0000 75.1500 160.6000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 160.0000 74.1500 160.6000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.0500 160.0000 73.1500 160.6000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.0500 160.0000 72.1500 160.6000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.0500 160.0000 71.1500 160.6000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.0500 160.0000 70.1500 160.6000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.0500 160.0000 69.1500 160.6000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.0500 160.0000 68.1500 160.6000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.0500 160.0000 67.1500 160.6000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.0500 160.0000 66.1500 160.6000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.0500 160.0000 65.1500 160.6000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.0500 160.0000 64.1500 160.6000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.0500 160.0000 63.1500 160.6000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.0500 160.0000 62.1500 160.6000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.0500 160.0000 61.1500 160.6000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.0500 160.0000 60.1500 160.6000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.0500 160.0000 59.1500 160.6000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.0500 160.0000 58.1500 160.6000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.0500 160.0000 57.1500 160.6000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.0500 160.0000 56.1500 160.6000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0500 160.0000 55.1500 160.6000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.0500 160.0000 54.1500 160.6000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.0500 160.0000 53.1500 160.6000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.0500 160.0000 52.1500 160.6000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.0500 160.0000 51.1500 160.6000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.0500 160.0000 50.1500 160.6000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.0500 160.0000 49.1500 160.6000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.0500 160.0000 48.1500 160.6000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.0500 160.0000 47.1500 160.6000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.0500 160.0000 46.1500 160.6000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.0500 160.0000 45.1500 160.6000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.0500 160.0000 44.1500 160.6000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.0500 160.0000 43.1500 160.6000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.0500 160.0000 42.1500 160.6000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.0500 160.0000 41.1500 160.6000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.0500 160.0000 40.1500 160.6000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.0500 160.0000 39.1500 160.6000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.0500 160.0000 38.1500 160.6000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.0500 160.0000 37.1500 160.6000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.0500 160.0000 36.1500 160.6000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.0500 160.0000 35.1500 160.6000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.0500 160.0000 34.1500 160.6000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0500 160.0000 33.1500 160.6000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.0500 160.0000 32.1500 160.6000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.0500 160.0000 31.1500 160.6000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.0500 160.0000 30.1500 160.6000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0500 160.0000 29.1500 160.6000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.0500 160.0000 28.1500 160.6000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.0500 160.0000 27.1500 160.6000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.0500 160.0000 26.1500 160.6000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.0500 160.0000 25.1500 160.6000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.0500 160.0000 24.1500 160.6000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.0500 160.0000 23.1500 160.6000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.0500 160.0000 22.1500 160.6000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.0500 160.0000 21.1500 160.6000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.0500 160.0000 20.1500 160.6000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.0500 160.0000 19.1500 160.6000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 160.0000 18.1500 160.6000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 76.3500 0.6000 76.4500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.3500 0.6000 72.4500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 80.3500 0.6000 80.4500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 84.3500 0.6000 84.4500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 88.3500 0.6000 88.4500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 92.3500 0.6000 92.4500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 12.0000 2.0000 14.0000 158.6000 ;
        RECT 28.2200 2.0000 30.2200 158.6000 ;
        RECT 44.4400 2.0000 46.4400 158.6000 ;
        RECT 60.6600 2.0000 62.6600 158.6000 ;
        RECT 76.8800 2.0000 78.8800 158.6000 ;
        RECT 93.1000 2.0000 95.1000 158.6000 ;
        RECT 109.3200 2.0000 111.3200 158.6000 ;
        RECT 125.5400 2.0000 127.5400 158.6000 ;
        RECT 141.7600 2.0000 143.7600 158.6000 ;
        RECT 157.9800 2.0000 159.9800 158.6000 ;
        RECT 12.0000 158.4350 14.0000 158.7650 ;
        RECT 28.2200 158.4350 30.2200 158.7650 ;
        RECT 60.6600 158.4350 62.6600 158.7650 ;
        RECT 44.4400 158.4350 46.4400 158.7650 ;
        RECT 76.8800 158.4350 78.8800 158.7650 ;
        RECT 93.1000 158.4350 95.1000 158.7650 ;
        RECT 109.3200 158.4350 111.3200 158.7650 ;
        RECT 141.7600 158.4350 143.7600 158.7650 ;
        RECT 125.5400 158.4350 127.5400 158.7650 ;
        RECT 157.9800 158.4350 159.9800 158.7650 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 5.0000 2.0000 7.0000 158.6000 ;
        RECT 21.2200 2.0000 23.2200 158.6000 ;
        RECT 37.4400 2.0000 39.4400 158.6000 ;
        RECT 53.6600 2.0000 55.6600 158.6000 ;
        RECT 69.8800 2.0000 71.8800 158.6000 ;
        RECT 86.1000 2.0000 88.1000 158.6000 ;
        RECT 102.3200 2.0000 104.3200 158.6000 ;
        RECT 118.5400 2.0000 120.5400 158.6000 ;
        RECT 134.7600 2.0000 136.7600 158.6000 ;
        RECT 150.9800 2.0000 152.9800 158.6000 ;
        RECT 5.0000 1.8350 7.0000 2.1650 ;
        RECT 21.2200 1.8350 23.2200 2.1650 ;
        RECT 37.4400 1.8350 39.4400 2.1650 ;
        RECT 53.6600 1.8350 55.6600 2.1650 ;
        RECT 69.8800 1.8350 71.8800 2.1650 ;
        RECT 102.3200 1.8350 104.3200 2.1650 ;
        RECT 86.1000 1.8350 88.1000 2.1650 ;
        RECT 118.5400 1.8350 120.5400 2.1650 ;
        RECT 134.7600 1.8350 136.7600 2.1650 ;
        RECT 150.9800 1.8350 152.9800 2.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 163.8000 160.6000 ;
    LAYER M2 ;
      RECT 145.2500 159.9000 163.8000 160.6000 ;
      RECT 144.2500 159.9000 144.9500 160.6000 ;
      RECT 143.2500 159.9000 143.9500 160.6000 ;
      RECT 142.2500 159.9000 142.9500 160.6000 ;
      RECT 141.2500 159.9000 141.9500 160.6000 ;
      RECT 140.2500 159.9000 140.9500 160.6000 ;
      RECT 139.2500 159.9000 139.9500 160.6000 ;
      RECT 138.2500 159.9000 138.9500 160.6000 ;
      RECT 137.2500 159.9000 137.9500 160.6000 ;
      RECT 136.2500 159.9000 136.9500 160.6000 ;
      RECT 135.2500 159.9000 135.9500 160.6000 ;
      RECT 134.2500 159.9000 134.9500 160.6000 ;
      RECT 133.2500 159.9000 133.9500 160.6000 ;
      RECT 132.2500 159.9000 132.9500 160.6000 ;
      RECT 131.2500 159.9000 131.9500 160.6000 ;
      RECT 130.2500 159.9000 130.9500 160.6000 ;
      RECT 129.2500 159.9000 129.9500 160.6000 ;
      RECT 128.2500 159.9000 128.9500 160.6000 ;
      RECT 127.2500 159.9000 127.9500 160.6000 ;
      RECT 126.2500 159.9000 126.9500 160.6000 ;
      RECT 125.2500 159.9000 125.9500 160.6000 ;
      RECT 124.2500 159.9000 124.9500 160.6000 ;
      RECT 123.2500 159.9000 123.9500 160.6000 ;
      RECT 122.2500 159.9000 122.9500 160.6000 ;
      RECT 121.2500 159.9000 121.9500 160.6000 ;
      RECT 120.2500 159.9000 120.9500 160.6000 ;
      RECT 119.2500 159.9000 119.9500 160.6000 ;
      RECT 118.2500 159.9000 118.9500 160.6000 ;
      RECT 117.2500 159.9000 117.9500 160.6000 ;
      RECT 116.2500 159.9000 116.9500 160.6000 ;
      RECT 115.2500 159.9000 115.9500 160.6000 ;
      RECT 114.2500 159.9000 114.9500 160.6000 ;
      RECT 113.2500 159.9000 113.9500 160.6000 ;
      RECT 112.2500 159.9000 112.9500 160.6000 ;
      RECT 111.2500 159.9000 111.9500 160.6000 ;
      RECT 110.2500 159.9000 110.9500 160.6000 ;
      RECT 109.2500 159.9000 109.9500 160.6000 ;
      RECT 108.2500 159.9000 108.9500 160.6000 ;
      RECT 107.2500 159.9000 107.9500 160.6000 ;
      RECT 106.2500 159.9000 106.9500 160.6000 ;
      RECT 105.2500 159.9000 105.9500 160.6000 ;
      RECT 104.2500 159.9000 104.9500 160.6000 ;
      RECT 103.2500 159.9000 103.9500 160.6000 ;
      RECT 102.2500 159.9000 102.9500 160.6000 ;
      RECT 101.2500 159.9000 101.9500 160.6000 ;
      RECT 100.2500 159.9000 100.9500 160.6000 ;
      RECT 99.2500 159.9000 99.9500 160.6000 ;
      RECT 98.2500 159.9000 98.9500 160.6000 ;
      RECT 97.2500 159.9000 97.9500 160.6000 ;
      RECT 96.2500 159.9000 96.9500 160.6000 ;
      RECT 95.2500 159.9000 95.9500 160.6000 ;
      RECT 94.2500 159.9000 94.9500 160.6000 ;
      RECT 93.2500 159.9000 93.9500 160.6000 ;
      RECT 92.2500 159.9000 92.9500 160.6000 ;
      RECT 91.2500 159.9000 91.9500 160.6000 ;
      RECT 90.2500 159.9000 90.9500 160.6000 ;
      RECT 89.2500 159.9000 89.9500 160.6000 ;
      RECT 88.2500 159.9000 88.9500 160.6000 ;
      RECT 87.2500 159.9000 87.9500 160.6000 ;
      RECT 86.2500 159.9000 86.9500 160.6000 ;
      RECT 85.2500 159.9000 85.9500 160.6000 ;
      RECT 84.2500 159.9000 84.9500 160.6000 ;
      RECT 83.2500 159.9000 83.9500 160.6000 ;
      RECT 82.2500 159.9000 82.9500 160.6000 ;
      RECT 81.2500 159.9000 81.9500 160.6000 ;
      RECT 80.2500 159.9000 80.9500 160.6000 ;
      RECT 79.2500 159.9000 79.9500 160.6000 ;
      RECT 78.2500 159.9000 78.9500 160.6000 ;
      RECT 77.2500 159.9000 77.9500 160.6000 ;
      RECT 76.2500 159.9000 76.9500 160.6000 ;
      RECT 75.2500 159.9000 75.9500 160.6000 ;
      RECT 74.2500 159.9000 74.9500 160.6000 ;
      RECT 73.2500 159.9000 73.9500 160.6000 ;
      RECT 72.2500 159.9000 72.9500 160.6000 ;
      RECT 71.2500 159.9000 71.9500 160.6000 ;
      RECT 70.2500 159.9000 70.9500 160.6000 ;
      RECT 69.2500 159.9000 69.9500 160.6000 ;
      RECT 68.2500 159.9000 68.9500 160.6000 ;
      RECT 67.2500 159.9000 67.9500 160.6000 ;
      RECT 66.2500 159.9000 66.9500 160.6000 ;
      RECT 65.2500 159.9000 65.9500 160.6000 ;
      RECT 64.2500 159.9000 64.9500 160.6000 ;
      RECT 63.2500 159.9000 63.9500 160.6000 ;
      RECT 62.2500 159.9000 62.9500 160.6000 ;
      RECT 61.2500 159.9000 61.9500 160.6000 ;
      RECT 60.2500 159.9000 60.9500 160.6000 ;
      RECT 59.2500 159.9000 59.9500 160.6000 ;
      RECT 58.2500 159.9000 58.9500 160.6000 ;
      RECT 57.2500 159.9000 57.9500 160.6000 ;
      RECT 56.2500 159.9000 56.9500 160.6000 ;
      RECT 55.2500 159.9000 55.9500 160.6000 ;
      RECT 54.2500 159.9000 54.9500 160.6000 ;
      RECT 53.2500 159.9000 53.9500 160.6000 ;
      RECT 52.2500 159.9000 52.9500 160.6000 ;
      RECT 51.2500 159.9000 51.9500 160.6000 ;
      RECT 50.2500 159.9000 50.9500 160.6000 ;
      RECT 49.2500 159.9000 49.9500 160.6000 ;
      RECT 48.2500 159.9000 48.9500 160.6000 ;
      RECT 47.2500 159.9000 47.9500 160.6000 ;
      RECT 46.2500 159.9000 46.9500 160.6000 ;
      RECT 45.2500 159.9000 45.9500 160.6000 ;
      RECT 44.2500 159.9000 44.9500 160.6000 ;
      RECT 43.2500 159.9000 43.9500 160.6000 ;
      RECT 42.2500 159.9000 42.9500 160.6000 ;
      RECT 41.2500 159.9000 41.9500 160.6000 ;
      RECT 40.2500 159.9000 40.9500 160.6000 ;
      RECT 39.2500 159.9000 39.9500 160.6000 ;
      RECT 38.2500 159.9000 38.9500 160.6000 ;
      RECT 37.2500 159.9000 37.9500 160.6000 ;
      RECT 36.2500 159.9000 36.9500 160.6000 ;
      RECT 35.2500 159.9000 35.9500 160.6000 ;
      RECT 34.2500 159.9000 34.9500 160.6000 ;
      RECT 33.2500 159.9000 33.9500 160.6000 ;
      RECT 32.2500 159.9000 32.9500 160.6000 ;
      RECT 31.2500 159.9000 31.9500 160.6000 ;
      RECT 30.2500 159.9000 30.9500 160.6000 ;
      RECT 29.2500 159.9000 29.9500 160.6000 ;
      RECT 28.2500 159.9000 28.9500 160.6000 ;
      RECT 27.2500 159.9000 27.9500 160.6000 ;
      RECT 26.2500 159.9000 26.9500 160.6000 ;
      RECT 25.2500 159.9000 25.9500 160.6000 ;
      RECT 24.2500 159.9000 24.9500 160.6000 ;
      RECT 23.2500 159.9000 23.9500 160.6000 ;
      RECT 22.2500 159.9000 22.9500 160.6000 ;
      RECT 21.2500 159.9000 21.9500 160.6000 ;
      RECT 20.2500 159.9000 20.9500 160.6000 ;
      RECT 19.2500 159.9000 19.9500 160.6000 ;
      RECT 18.2500 159.9000 18.9500 160.6000 ;
      RECT 0.0000 159.9000 17.9500 160.6000 ;
      RECT 0.0000 0.7000 163.8000 159.9000 ;
      RECT 145.2500 0.0000 163.8000 0.7000 ;
      RECT 144.2500 0.0000 144.9500 0.7000 ;
      RECT 143.2500 0.0000 143.9500 0.7000 ;
      RECT 142.2500 0.0000 142.9500 0.7000 ;
      RECT 141.2500 0.0000 141.9500 0.7000 ;
      RECT 140.2500 0.0000 140.9500 0.7000 ;
      RECT 139.2500 0.0000 139.9500 0.7000 ;
      RECT 138.2500 0.0000 138.9500 0.7000 ;
      RECT 137.2500 0.0000 137.9500 0.7000 ;
      RECT 136.2500 0.0000 136.9500 0.7000 ;
      RECT 135.2500 0.0000 135.9500 0.7000 ;
      RECT 134.2500 0.0000 134.9500 0.7000 ;
      RECT 133.2500 0.0000 133.9500 0.7000 ;
      RECT 132.2500 0.0000 132.9500 0.7000 ;
      RECT 131.2500 0.0000 131.9500 0.7000 ;
      RECT 130.2500 0.0000 130.9500 0.7000 ;
      RECT 129.2500 0.0000 129.9500 0.7000 ;
      RECT 128.2500 0.0000 128.9500 0.7000 ;
      RECT 127.2500 0.0000 127.9500 0.7000 ;
      RECT 126.2500 0.0000 126.9500 0.7000 ;
      RECT 125.2500 0.0000 125.9500 0.7000 ;
      RECT 124.2500 0.0000 124.9500 0.7000 ;
      RECT 123.2500 0.0000 123.9500 0.7000 ;
      RECT 122.2500 0.0000 122.9500 0.7000 ;
      RECT 121.2500 0.0000 121.9500 0.7000 ;
      RECT 120.2500 0.0000 120.9500 0.7000 ;
      RECT 119.2500 0.0000 119.9500 0.7000 ;
      RECT 118.2500 0.0000 118.9500 0.7000 ;
      RECT 117.2500 0.0000 117.9500 0.7000 ;
      RECT 116.2500 0.0000 116.9500 0.7000 ;
      RECT 115.2500 0.0000 115.9500 0.7000 ;
      RECT 114.2500 0.0000 114.9500 0.7000 ;
      RECT 113.2500 0.0000 113.9500 0.7000 ;
      RECT 112.2500 0.0000 112.9500 0.7000 ;
      RECT 111.2500 0.0000 111.9500 0.7000 ;
      RECT 110.2500 0.0000 110.9500 0.7000 ;
      RECT 109.2500 0.0000 109.9500 0.7000 ;
      RECT 108.2500 0.0000 108.9500 0.7000 ;
      RECT 107.2500 0.0000 107.9500 0.7000 ;
      RECT 106.2500 0.0000 106.9500 0.7000 ;
      RECT 105.2500 0.0000 105.9500 0.7000 ;
      RECT 104.2500 0.0000 104.9500 0.7000 ;
      RECT 103.2500 0.0000 103.9500 0.7000 ;
      RECT 102.2500 0.0000 102.9500 0.7000 ;
      RECT 101.2500 0.0000 101.9500 0.7000 ;
      RECT 100.2500 0.0000 100.9500 0.7000 ;
      RECT 99.2500 0.0000 99.9500 0.7000 ;
      RECT 98.2500 0.0000 98.9500 0.7000 ;
      RECT 97.2500 0.0000 97.9500 0.7000 ;
      RECT 96.2500 0.0000 96.9500 0.7000 ;
      RECT 95.2500 0.0000 95.9500 0.7000 ;
      RECT 94.2500 0.0000 94.9500 0.7000 ;
      RECT 93.2500 0.0000 93.9500 0.7000 ;
      RECT 92.2500 0.0000 92.9500 0.7000 ;
      RECT 91.2500 0.0000 91.9500 0.7000 ;
      RECT 90.2500 0.0000 90.9500 0.7000 ;
      RECT 89.2500 0.0000 89.9500 0.7000 ;
      RECT 88.2500 0.0000 88.9500 0.7000 ;
      RECT 87.2500 0.0000 87.9500 0.7000 ;
      RECT 86.2500 0.0000 86.9500 0.7000 ;
      RECT 85.2500 0.0000 85.9500 0.7000 ;
      RECT 84.2500 0.0000 84.9500 0.7000 ;
      RECT 83.2500 0.0000 83.9500 0.7000 ;
      RECT 82.2500 0.0000 82.9500 0.7000 ;
      RECT 81.2500 0.0000 81.9500 0.7000 ;
      RECT 80.2500 0.0000 80.9500 0.7000 ;
      RECT 79.2500 0.0000 79.9500 0.7000 ;
      RECT 78.2500 0.0000 78.9500 0.7000 ;
      RECT 77.2500 0.0000 77.9500 0.7000 ;
      RECT 76.2500 0.0000 76.9500 0.7000 ;
      RECT 75.2500 0.0000 75.9500 0.7000 ;
      RECT 74.2500 0.0000 74.9500 0.7000 ;
      RECT 73.2500 0.0000 73.9500 0.7000 ;
      RECT 72.2500 0.0000 72.9500 0.7000 ;
      RECT 71.2500 0.0000 71.9500 0.7000 ;
      RECT 70.2500 0.0000 70.9500 0.7000 ;
      RECT 69.2500 0.0000 69.9500 0.7000 ;
      RECT 68.2500 0.0000 68.9500 0.7000 ;
      RECT 67.2500 0.0000 67.9500 0.7000 ;
      RECT 66.2500 0.0000 66.9500 0.7000 ;
      RECT 65.2500 0.0000 65.9500 0.7000 ;
      RECT 64.2500 0.0000 64.9500 0.7000 ;
      RECT 63.2500 0.0000 63.9500 0.7000 ;
      RECT 62.2500 0.0000 62.9500 0.7000 ;
      RECT 61.2500 0.0000 61.9500 0.7000 ;
      RECT 60.2500 0.0000 60.9500 0.7000 ;
      RECT 59.2500 0.0000 59.9500 0.7000 ;
      RECT 58.2500 0.0000 58.9500 0.7000 ;
      RECT 57.2500 0.0000 57.9500 0.7000 ;
      RECT 56.2500 0.0000 56.9500 0.7000 ;
      RECT 55.2500 0.0000 55.9500 0.7000 ;
      RECT 54.2500 0.0000 54.9500 0.7000 ;
      RECT 53.2500 0.0000 53.9500 0.7000 ;
      RECT 52.2500 0.0000 52.9500 0.7000 ;
      RECT 51.2500 0.0000 51.9500 0.7000 ;
      RECT 50.2500 0.0000 50.9500 0.7000 ;
      RECT 49.2500 0.0000 49.9500 0.7000 ;
      RECT 48.2500 0.0000 48.9500 0.7000 ;
      RECT 47.2500 0.0000 47.9500 0.7000 ;
      RECT 46.2500 0.0000 46.9500 0.7000 ;
      RECT 45.2500 0.0000 45.9500 0.7000 ;
      RECT 44.2500 0.0000 44.9500 0.7000 ;
      RECT 43.2500 0.0000 43.9500 0.7000 ;
      RECT 42.2500 0.0000 42.9500 0.7000 ;
      RECT 41.2500 0.0000 41.9500 0.7000 ;
      RECT 40.2500 0.0000 40.9500 0.7000 ;
      RECT 39.2500 0.0000 39.9500 0.7000 ;
      RECT 38.2500 0.0000 38.9500 0.7000 ;
      RECT 37.2500 0.0000 37.9500 0.7000 ;
      RECT 36.2500 0.0000 36.9500 0.7000 ;
      RECT 35.2500 0.0000 35.9500 0.7000 ;
      RECT 34.2500 0.0000 34.9500 0.7000 ;
      RECT 33.2500 0.0000 33.9500 0.7000 ;
      RECT 32.2500 0.0000 32.9500 0.7000 ;
      RECT 31.2500 0.0000 31.9500 0.7000 ;
      RECT 30.2500 0.0000 30.9500 0.7000 ;
      RECT 29.2500 0.0000 29.9500 0.7000 ;
      RECT 28.2500 0.0000 28.9500 0.7000 ;
      RECT 27.2500 0.0000 27.9500 0.7000 ;
      RECT 26.2500 0.0000 26.9500 0.7000 ;
      RECT 25.2500 0.0000 25.9500 0.7000 ;
      RECT 24.2500 0.0000 24.9500 0.7000 ;
      RECT 23.2500 0.0000 23.9500 0.7000 ;
      RECT 22.2500 0.0000 22.9500 0.7000 ;
      RECT 21.2500 0.0000 21.9500 0.7000 ;
      RECT 20.2500 0.0000 20.9500 0.7000 ;
      RECT 19.2500 0.0000 19.9500 0.7000 ;
      RECT 18.2500 0.0000 18.9500 0.7000 ;
      RECT 0.0000 0.0000 17.9500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 92.5500 163.8000 160.6000 ;
      RECT 0.7000 92.2500 163.8000 92.5500 ;
      RECT 0.0000 88.5500 163.8000 92.2500 ;
      RECT 0.7000 88.2500 163.8000 88.5500 ;
      RECT 0.0000 84.5500 163.8000 88.2500 ;
      RECT 0.7000 84.2500 163.8000 84.5500 ;
      RECT 0.0000 80.5500 163.8000 84.2500 ;
      RECT 0.7000 80.2500 163.8000 80.5500 ;
      RECT 0.0000 76.5500 163.8000 80.2500 ;
      RECT 0.7000 76.2500 163.8000 76.5500 ;
      RECT 0.0000 72.5500 163.8000 76.2500 ;
      RECT 0.7000 72.2500 163.8000 72.5500 ;
      RECT 0.0000 68.5500 163.8000 72.2500 ;
      RECT 0.7000 68.2500 163.8000 68.5500 ;
      RECT 0.0000 0.0000 163.8000 68.2500 ;
    LAYER M4 ;
      RECT 0.0000 159.2650 163.8000 160.6000 ;
      RECT 144.2600 159.1000 157.4800 159.2650 ;
      RECT 128.0400 159.1000 141.2600 159.2650 ;
      RECT 111.8200 159.1000 125.0400 159.2650 ;
      RECT 95.6000 159.1000 108.8200 159.2650 ;
      RECT 79.3800 159.1000 92.6000 159.2650 ;
      RECT 63.1600 159.1000 76.3800 159.2650 ;
      RECT 46.9400 159.1000 60.1600 159.2650 ;
      RECT 30.7200 159.1000 43.9400 159.2650 ;
      RECT 14.5000 159.1000 27.7200 159.2650 ;
      RECT 0.0000 159.1000 11.5000 159.2650 ;
      RECT 160.4800 1.5000 163.8000 159.2650 ;
      RECT 153.4800 1.5000 157.4800 159.1000 ;
      RECT 144.2600 1.5000 150.4800 159.1000 ;
      RECT 137.2600 1.5000 141.2600 159.1000 ;
      RECT 128.0400 1.5000 134.2600 159.1000 ;
      RECT 121.0400 1.5000 125.0400 159.1000 ;
      RECT 111.8200 1.5000 118.0400 159.1000 ;
      RECT 104.8200 1.5000 108.8200 159.1000 ;
      RECT 95.6000 1.5000 101.8200 159.1000 ;
      RECT 88.6000 1.5000 92.6000 159.1000 ;
      RECT 79.3800 1.5000 85.6000 159.1000 ;
      RECT 72.3800 1.5000 76.3800 159.1000 ;
      RECT 63.1600 1.5000 69.3800 159.1000 ;
      RECT 56.1600 1.5000 60.1600 159.1000 ;
      RECT 46.9400 1.5000 53.1600 159.1000 ;
      RECT 39.9400 1.5000 43.9400 159.1000 ;
      RECT 30.7200 1.5000 36.9400 159.1000 ;
      RECT 23.7200 1.5000 27.7200 159.1000 ;
      RECT 14.5000 1.5000 20.7200 159.1000 ;
      RECT 7.5000 1.5000 11.5000 159.1000 ;
      RECT 153.4800 1.3350 163.8000 1.5000 ;
      RECT 137.2600 1.3350 150.4800 1.5000 ;
      RECT 121.0400 1.3350 134.2600 1.5000 ;
      RECT 104.8200 1.3350 118.0400 1.5000 ;
      RECT 88.6000 1.3350 101.8200 1.5000 ;
      RECT 72.3800 1.3350 85.6000 1.5000 ;
      RECT 56.1600 1.3350 69.3800 1.5000 ;
      RECT 39.9400 1.3350 53.1600 1.5000 ;
      RECT 23.7200 1.3350 36.9400 1.5000 ;
      RECT 7.5000 1.3350 20.7200 1.5000 ;
      RECT 0.0000 1.3350 4.5000 159.1000 ;
      RECT 0.0000 0.0000 163.8000 1.3350 ;
  END
END sram_w8

END LIBRARY
