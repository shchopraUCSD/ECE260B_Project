##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 21:12:07 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 1761.4000 BY 1760.6000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 668.9500 0.5200 669.0500 ;
    END
  END clk1
  PIN clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 668.9500 1761.4000 669.0500 ;
    END
  END clk2
  PIN mem_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 664.9500 1761.4000 665.0500 ;
    END
  END mem_in[127]
  PIN mem_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 660.9500 1761.4000 661.0500 ;
    END
  END mem_in[126]
  PIN mem_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 656.9500 1761.4000 657.0500 ;
    END
  END mem_in[125]
  PIN mem_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 652.9500 1761.4000 653.0500 ;
    END
  END mem_in[124]
  PIN mem_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 648.9500 1761.4000 649.0500 ;
    END
  END mem_in[123]
  PIN mem_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 644.9500 1761.4000 645.0500 ;
    END
  END mem_in[122]
  PIN mem_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 640.9500 1761.4000 641.0500 ;
    END
  END mem_in[121]
  PIN mem_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 636.9500 1761.4000 637.0500 ;
    END
  END mem_in[120]
  PIN mem_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 632.9500 1761.4000 633.0500 ;
    END
  END mem_in[119]
  PIN mem_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 628.9500 1761.4000 629.0500 ;
    END
  END mem_in[118]
  PIN mem_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 624.9500 1761.4000 625.0500 ;
    END
  END mem_in[117]
  PIN mem_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 620.9500 1761.4000 621.0500 ;
    END
  END mem_in[116]
  PIN mem_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 616.9500 1761.4000 617.0500 ;
    END
  END mem_in[115]
  PIN mem_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 612.9500 1761.4000 613.0500 ;
    END
  END mem_in[114]
  PIN mem_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 608.9500 1761.4000 609.0500 ;
    END
  END mem_in[113]
  PIN mem_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 604.9500 1761.4000 605.0500 ;
    END
  END mem_in[112]
  PIN mem_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 600.9500 1761.4000 601.0500 ;
    END
  END mem_in[111]
  PIN mem_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 596.9500 1761.4000 597.0500 ;
    END
  END mem_in[110]
  PIN mem_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 592.9500 1761.4000 593.0500 ;
    END
  END mem_in[109]
  PIN mem_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 588.9500 1761.4000 589.0500 ;
    END
  END mem_in[108]
  PIN mem_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 584.9500 1761.4000 585.0500 ;
    END
  END mem_in[107]
  PIN mem_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 580.9500 1761.4000 581.0500 ;
    END
  END mem_in[106]
  PIN mem_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 576.9500 1761.4000 577.0500 ;
    END
  END mem_in[105]
  PIN mem_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 572.9500 1761.4000 573.0500 ;
    END
  END mem_in[104]
  PIN mem_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 568.9500 1761.4000 569.0500 ;
    END
  END mem_in[103]
  PIN mem_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 564.9500 1761.4000 565.0500 ;
    END
  END mem_in[102]
  PIN mem_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 560.9500 1761.4000 561.0500 ;
    END
  END mem_in[101]
  PIN mem_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 556.9500 1761.4000 557.0500 ;
    END
  END mem_in[100]
  PIN mem_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 552.9500 1761.4000 553.0500 ;
    END
  END mem_in[99]
  PIN mem_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 548.9500 1761.4000 549.0500 ;
    END
  END mem_in[98]
  PIN mem_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 544.9500 1761.4000 545.0500 ;
    END
  END mem_in[97]
  PIN mem_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 540.9500 1761.4000 541.0500 ;
    END
  END mem_in[96]
  PIN mem_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 536.9500 1761.4000 537.0500 ;
    END
  END mem_in[95]
  PIN mem_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 532.9500 1761.4000 533.0500 ;
    END
  END mem_in[94]
  PIN mem_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 528.9500 1761.4000 529.0500 ;
    END
  END mem_in[93]
  PIN mem_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 524.9500 1761.4000 525.0500 ;
    END
  END mem_in[92]
  PIN mem_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 520.9500 1761.4000 521.0500 ;
    END
  END mem_in[91]
  PIN mem_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 516.9500 1761.4000 517.0500 ;
    END
  END mem_in[90]
  PIN mem_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 512.9500 1761.4000 513.0500 ;
    END
  END mem_in[89]
  PIN mem_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 508.9500 1761.4000 509.0500 ;
    END
  END mem_in[88]
  PIN mem_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 504.9500 1761.4000 505.0500 ;
    END
  END mem_in[87]
  PIN mem_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 500.9500 1761.4000 501.0500 ;
    END
  END mem_in[86]
  PIN mem_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 496.9500 1761.4000 497.0500 ;
    END
  END mem_in[85]
  PIN mem_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 492.9500 1761.4000 493.0500 ;
    END
  END mem_in[84]
  PIN mem_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 488.9500 1761.4000 489.0500 ;
    END
  END mem_in[83]
  PIN mem_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 484.9500 1761.4000 485.0500 ;
    END
  END mem_in[82]
  PIN mem_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 480.9500 1761.4000 481.0500 ;
    END
  END mem_in[81]
  PIN mem_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 476.9500 1761.4000 477.0500 ;
    END
  END mem_in[80]
  PIN mem_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 472.9500 1761.4000 473.0500 ;
    END
  END mem_in[79]
  PIN mem_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 468.9500 1761.4000 469.0500 ;
    END
  END mem_in[78]
  PIN mem_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 464.9500 1761.4000 465.0500 ;
    END
  END mem_in[77]
  PIN mem_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 460.9500 1761.4000 461.0500 ;
    END
  END mem_in[76]
  PIN mem_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 456.9500 1761.4000 457.0500 ;
    END
  END mem_in[75]
  PIN mem_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 452.9500 1761.4000 453.0500 ;
    END
  END mem_in[74]
  PIN mem_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 448.9500 1761.4000 449.0500 ;
    END
  END mem_in[73]
  PIN mem_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 444.9500 1761.4000 445.0500 ;
    END
  END mem_in[72]
  PIN mem_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 440.9500 1761.4000 441.0500 ;
    END
  END mem_in[71]
  PIN mem_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 436.9500 1761.4000 437.0500 ;
    END
  END mem_in[70]
  PIN mem_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 432.9500 1761.4000 433.0500 ;
    END
  END mem_in[69]
  PIN mem_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 428.9500 1761.4000 429.0500 ;
    END
  END mem_in[68]
  PIN mem_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 424.9500 1761.4000 425.0500 ;
    END
  END mem_in[67]
  PIN mem_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 420.9500 1761.4000 421.0500 ;
    END
  END mem_in[66]
  PIN mem_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 416.9500 1761.4000 417.0500 ;
    END
  END mem_in[65]
  PIN mem_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 412.9500 1761.4000 413.0500 ;
    END
  END mem_in[64]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 664.9500 0.5200 665.0500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 660.9500 0.5200 661.0500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 656.9500 0.5200 657.0500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 652.9500 0.5200 653.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 648.9500 0.5200 649.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 644.9500 0.5200 645.0500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 640.9500 0.5200 641.0500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 636.9500 0.5200 637.0500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 632.9500 0.5200 633.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 628.9500 0.5200 629.0500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 624.9500 0.5200 625.0500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 620.9500 0.5200 621.0500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 616.9500 0.5200 617.0500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 612.9500 0.5200 613.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 608.9500 0.5200 609.0500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 604.9500 0.5200 605.0500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 600.9500 0.5200 601.0500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 596.9500 0.5200 597.0500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 592.9500 0.5200 593.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 588.9500 0.5200 589.0500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 584.9500 0.5200 585.0500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 580.9500 0.5200 581.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 576.9500 0.5200 577.0500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 572.9500 0.5200 573.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 568.9500 0.5200 569.0500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 564.9500 0.5200 565.0500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 560.9500 0.5200 561.0500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 556.9500 0.5200 557.0500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 552.9500 0.5200 553.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 548.9500 0.5200 549.0500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 544.9500 0.5200 545.0500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 540.9500 0.5200 541.0500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 536.9500 0.5200 537.0500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 532.9500 0.5200 533.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 528.9500 0.5200 529.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 524.9500 0.5200 525.0500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 520.9500 0.5200 521.0500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 516.9500 0.5200 517.0500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 512.9500 0.5200 513.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 508.9500 0.5200 509.0500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 504.9500 0.5200 505.0500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 500.9500 0.5200 501.0500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 496.9500 0.5200 497.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 492.9500 0.5200 493.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 488.9500 0.5200 489.0500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 484.9500 0.5200 485.0500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 480.9500 0.5200 481.0500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 476.9500 0.5200 477.0500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 472.9500 0.5200 473.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 468.9500 0.5200 469.0500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 464.9500 0.5200 465.0500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 460.9500 0.5200 461.0500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 456.9500 0.5200 457.0500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 452.9500 0.5200 453.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 448.9500 0.5200 449.0500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 444.9500 0.5200 445.0500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 440.9500 0.5200 441.0500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 436.9500 0.5200 437.0500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 432.9500 0.5200 433.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 428.9500 0.5200 429.0500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 424.9500 0.5200 425.0500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 420.9500 0.5200 421.0500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 416.9500 0.5200 417.0500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 412.9500 0.5200 413.0500 ;
    END
  END mem_in[0]
  PIN inst[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 408.9500 1761.4000 409.0500 ;
    END
  END inst[43]
  PIN inst[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 404.9500 1761.4000 405.0500 ;
    END
  END inst[42]
  PIN inst[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 400.9500 1761.4000 401.0500 ;
    END
  END inst[41]
  PIN inst[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 396.9500 1761.4000 397.0500 ;
    END
  END inst[40]
  PIN inst[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 392.9500 1761.4000 393.0500 ;
    END
  END inst[39]
  PIN inst[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 388.9500 1761.4000 389.0500 ;
    END
  END inst[38]
  PIN inst[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 384.9500 1761.4000 385.0500 ;
    END
  END inst[37]
  PIN inst[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 380.9500 1761.4000 381.0500 ;
    END
  END inst[36]
  PIN inst[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 376.9500 1761.4000 377.0500 ;
    END
  END inst[35]
  PIN inst[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 372.9500 1761.4000 373.0500 ;
    END
  END inst[34]
  PIN inst[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 368.9500 1761.4000 369.0500 ;
    END
  END inst[33]
  PIN inst[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 364.9500 1761.4000 365.0500 ;
    END
  END inst[32]
  PIN inst[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 360.9500 1761.4000 361.0500 ;
    END
  END inst[31]
  PIN inst[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 356.9500 1761.4000 357.0500 ;
    END
  END inst[30]
  PIN inst[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 352.9500 1761.4000 353.0500 ;
    END
  END inst[29]
  PIN inst[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 348.9500 1761.4000 349.0500 ;
    END
  END inst[28]
  PIN inst[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 344.9500 1761.4000 345.0500 ;
    END
  END inst[27]
  PIN inst[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 340.9500 1761.4000 341.0500 ;
    END
  END inst[26]
  PIN inst[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 336.9500 1761.4000 337.0500 ;
    END
  END inst[25]
  PIN inst[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 332.9500 1761.4000 333.0500 ;
    END
  END inst[24]
  PIN inst[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 328.9500 1761.4000 329.0500 ;
    END
  END inst[23]
  PIN inst[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1760.8800 324.9500 1761.4000 325.0500 ;
    END
  END inst[22]
  PIN inst[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 408.9500 0.5200 409.0500 ;
    END
  END inst[21]
  PIN inst[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 404.9500 0.5200 405.0500 ;
    END
  END inst[20]
  PIN inst[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 400.9500 0.5200 401.0500 ;
    END
  END inst[19]
  PIN inst[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 396.9500 0.5200 397.0500 ;
    END
  END inst[18]
  PIN inst[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 392.9500 0.5200 393.0500 ;
    END
  END inst[17]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 388.9500 0.5200 389.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 384.9500 0.5200 385.0500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 380.9500 0.5200 381.0500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 376.9500 0.5200 377.0500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 372.9500 0.5200 373.0500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 368.9500 0.5200 369.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 364.9500 0.5200 365.0500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 360.9500 0.5200 361.0500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 356.9500 0.5200 357.0500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 352.9500 0.5200 353.0500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 348.9500 0.5200 349.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 344.9500 0.5200 345.0500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 340.9500 0.5200 341.0500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 336.9500 0.5200 337.0500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 332.9500 0.5200 333.0500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 328.9500 0.5200 329.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 0.0000 324.9500 0.5200 325.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 880.8500 0.0000 880.9500 0.5200 ;
    END
  END reset
  PIN out[319]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1009.4500 0.0000 1009.5500 0.5200 ;
    END
  END out[319]
  PIN out[318]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1016.4500 0.0000 1016.5500 0.5200 ;
    END
  END out[318]
  PIN out[317]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1023.4500 0.0000 1023.5500 0.5200 ;
    END
  END out[317]
  PIN out[316]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1030.4500 0.0000 1030.5500 0.5200 ;
    END
  END out[316]
  PIN out[315]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1037.4500 0.0000 1037.5500 0.5200 ;
    END
  END out[315]
  PIN out[314]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1044.4500 0.0000 1044.5500 0.5200 ;
    END
  END out[314]
  PIN out[313]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1051.4500 0.0000 1051.5500 0.5200 ;
    END
  END out[313]
  PIN out[312]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1058.4500 0.0000 1058.5500 0.5200 ;
    END
  END out[312]
  PIN out[311]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1065.4500 0.0000 1065.5500 0.5200 ;
    END
  END out[311]
  PIN out[310]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1072.4500 0.0000 1072.5500 0.5200 ;
    END
  END out[310]
  PIN out[309]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1079.4500 0.0000 1079.5500 0.5200 ;
    END
  END out[309]
  PIN out[308]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1086.4500 0.0000 1086.5500 0.5200 ;
    END
  END out[308]
  PIN out[307]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1093.4500 0.0000 1093.5500 0.5200 ;
    END
  END out[307]
  PIN out[306]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1100.4500 0.0000 1100.5500 0.5200 ;
    END
  END out[306]
  PIN out[305]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1107.4500 0.0000 1107.5500 0.5200 ;
    END
  END out[305]
  PIN out[304]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1114.4500 0.0000 1114.5500 0.5200 ;
    END
  END out[304]
  PIN out[303]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1121.4500 0.0000 1121.5500 0.5200 ;
    END
  END out[303]
  PIN out[302]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1128.4500 0.0000 1128.5500 0.5200 ;
    END
  END out[302]
  PIN out[301]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1135.4500 0.0000 1135.5500 0.5200 ;
    END
  END out[301]
  PIN out[300]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1142.4500 0.0000 1142.5500 0.5200 ;
    END
  END out[300]
  PIN out[299]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1149.4500 0.0000 1149.5500 0.5200 ;
    END
  END out[299]
  PIN out[298]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1156.4500 0.0000 1156.5500 0.5200 ;
    END
  END out[298]
  PIN out[297]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1163.4500 0.0000 1163.5500 0.5200 ;
    END
  END out[297]
  PIN out[296]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1170.4500 0.0000 1170.5500 0.5200 ;
    END
  END out[296]
  PIN out[295]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1177.4500 0.0000 1177.5500 0.5200 ;
    END
  END out[295]
  PIN out[294]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1184.4500 0.0000 1184.5500 0.5200 ;
    END
  END out[294]
  PIN out[293]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1191.4500 0.0000 1191.5500 0.5200 ;
    END
  END out[293]
  PIN out[292]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1198.4500 0.0000 1198.5500 0.5200 ;
    END
  END out[292]
  PIN out[291]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1205.4500 0.0000 1205.5500 0.5200 ;
    END
  END out[291]
  PIN out[290]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1212.4500 0.0000 1212.5500 0.5200 ;
    END
  END out[290]
  PIN out[289]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1219.4500 0.0000 1219.5500 0.5200 ;
    END
  END out[289]
  PIN out[288]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1226.4500 0.0000 1226.5500 0.5200 ;
    END
  END out[288]
  PIN out[287]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1233.4500 0.0000 1233.5500 0.5200 ;
    END
  END out[287]
  PIN out[286]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1240.4500 0.0000 1240.5500 0.5200 ;
    END
  END out[286]
  PIN out[285]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1247.4500 0.0000 1247.5500 0.5200 ;
    END
  END out[285]
  PIN out[284]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1254.4500 0.0000 1254.5500 0.5200 ;
    END
  END out[284]
  PIN out[283]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1261.4500 0.0000 1261.5500 0.5200 ;
    END
  END out[283]
  PIN out[282]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1268.4500 0.0000 1268.5500 0.5200 ;
    END
  END out[282]
  PIN out[281]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1275.4500 0.0000 1275.5500 0.5200 ;
    END
  END out[281]
  PIN out[280]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1282.4500 0.0000 1282.5500 0.5200 ;
    END
  END out[280]
  PIN out[279]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1289.4500 0.0000 1289.5500 0.5200 ;
    END
  END out[279]
  PIN out[278]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1296.4500 0.0000 1296.5500 0.5200 ;
    END
  END out[278]
  PIN out[277]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1303.4500 0.0000 1303.5500 0.5200 ;
    END
  END out[277]
  PIN out[276]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1310.4500 0.0000 1310.5500 0.5200 ;
    END
  END out[276]
  PIN out[275]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1317.4500 0.0000 1317.5500 0.5200 ;
    END
  END out[275]
  PIN out[274]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1324.4500 0.0000 1324.5500 0.5200 ;
    END
  END out[274]
  PIN out[273]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1331.4500 0.0000 1331.5500 0.5200 ;
    END
  END out[273]
  PIN out[272]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1338.4500 0.0000 1338.5500 0.5200 ;
    END
  END out[272]
  PIN out[271]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1345.4500 0.0000 1345.5500 0.5200 ;
    END
  END out[271]
  PIN out[270]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1352.4500 0.0000 1352.5500 0.5200 ;
    END
  END out[270]
  PIN out[269]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1359.4500 0.0000 1359.5500 0.5200 ;
    END
  END out[269]
  PIN out[268]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1366.4500 0.0000 1366.5500 0.5200 ;
    END
  END out[268]
  PIN out[267]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1373.4500 0.0000 1373.5500 0.5200 ;
    END
  END out[267]
  PIN out[266]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1380.4500 0.0000 1380.5500 0.5200 ;
    END
  END out[266]
  PIN out[265]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1387.4500 0.0000 1387.5500 0.5200 ;
    END
  END out[265]
  PIN out[264]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1394.4500 0.0000 1394.5500 0.5200 ;
    END
  END out[264]
  PIN out[263]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1401.4500 0.0000 1401.5500 0.5200 ;
    END
  END out[263]
  PIN out[262]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1408.4500 0.0000 1408.5500 0.5200 ;
    END
  END out[262]
  PIN out[261]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1415.4500 0.0000 1415.5500 0.5200 ;
    END
  END out[261]
  PIN out[260]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1422.4500 0.0000 1422.5500 0.5200 ;
    END
  END out[260]
  PIN out[259]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1429.4500 0.0000 1429.5500 0.5200 ;
    END
  END out[259]
  PIN out[258]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1436.4500 0.0000 1436.5500 0.5200 ;
    END
  END out[258]
  PIN out[257]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1443.4500 0.0000 1443.5500 0.5200 ;
    END
  END out[257]
  PIN out[256]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1450.4500 0.0000 1450.5500 0.5200 ;
    END
  END out[256]
  PIN out[255]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1457.4500 0.0000 1457.5500 0.5200 ;
    END
  END out[255]
  PIN out[254]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1464.4500 0.0000 1464.5500 0.5200 ;
    END
  END out[254]
  PIN out[253]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1471.4500 0.0000 1471.5500 0.5200 ;
    END
  END out[253]
  PIN out[252]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1478.4500 0.0000 1478.5500 0.5200 ;
    END
  END out[252]
  PIN out[251]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1485.4500 0.0000 1485.5500 0.5200 ;
    END
  END out[251]
  PIN out[250]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1492.4500 0.0000 1492.5500 0.5200 ;
    END
  END out[250]
  PIN out[249]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1499.4500 0.0000 1499.5500 0.5200 ;
    END
  END out[249]
  PIN out[248]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1506.4500 0.0000 1506.5500 0.5200 ;
    END
  END out[248]
  PIN out[247]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1513.4500 0.0000 1513.5500 0.5200 ;
    END
  END out[247]
  PIN out[246]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1520.4500 0.0000 1520.5500 0.5200 ;
    END
  END out[246]
  PIN out[245]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1527.4500 0.0000 1527.5500 0.5200 ;
    END
  END out[245]
  PIN out[244]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1534.4500 0.0000 1534.5500 0.5200 ;
    END
  END out[244]
  PIN out[243]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1541.4500 0.0000 1541.5500 0.5200 ;
    END
  END out[243]
  PIN out[242]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1548.4500 0.0000 1548.5500 0.5200 ;
    END
  END out[242]
  PIN out[241]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1555.4500 0.0000 1555.5500 0.5200 ;
    END
  END out[241]
  PIN out[240]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1562.4500 0.0000 1562.5500 0.5200 ;
    END
  END out[240]
  PIN out[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1012.8500 0.0000 1012.9500 0.5200 ;
    END
  END out[239]
  PIN out[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1019.8500 0.0000 1019.9500 0.5200 ;
    END
  END out[238]
  PIN out[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1026.8500 0.0000 1026.9500 0.5200 ;
    END
  END out[237]
  PIN out[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1033.8500 0.0000 1033.9500 0.5200 ;
    END
  END out[236]
  PIN out[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1040.8500 0.0000 1040.9500 0.5200 ;
    END
  END out[235]
  PIN out[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1047.8500 0.0000 1047.9500 0.5200 ;
    END
  END out[234]
  PIN out[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1054.8500 0.0000 1054.9500 0.5200 ;
    END
  END out[233]
  PIN out[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1061.8500 0.0000 1061.9500 0.5200 ;
    END
  END out[232]
  PIN out[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1068.8500 0.0000 1068.9500 0.5200 ;
    END
  END out[231]
  PIN out[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1075.8500 0.0000 1075.9500 0.5200 ;
    END
  END out[230]
  PIN out[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1082.8500 0.0000 1082.9500 0.5200 ;
    END
  END out[229]
  PIN out[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1089.8500 0.0000 1089.9500 0.5200 ;
    END
  END out[228]
  PIN out[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1096.8500 0.0000 1096.9500 0.5200 ;
    END
  END out[227]
  PIN out[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1103.8500 0.0000 1103.9500 0.5200 ;
    END
  END out[226]
  PIN out[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1110.8500 0.0000 1110.9500 0.5200 ;
    END
  END out[225]
  PIN out[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1117.8500 0.0000 1117.9500 0.5200 ;
    END
  END out[224]
  PIN out[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1124.8500 0.0000 1124.9500 0.5200 ;
    END
  END out[223]
  PIN out[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1131.8500 0.0000 1131.9500 0.5200 ;
    END
  END out[222]
  PIN out[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1138.8500 0.0000 1138.9500 0.5200 ;
    END
  END out[221]
  PIN out[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1145.8500 0.0000 1145.9500 0.5200 ;
    END
  END out[220]
  PIN out[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1152.8500 0.0000 1152.9500 0.5200 ;
    END
  END out[219]
  PIN out[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1159.8500 0.0000 1159.9500 0.5200 ;
    END
  END out[218]
  PIN out[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1166.8500 0.0000 1166.9500 0.5200 ;
    END
  END out[217]
  PIN out[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1173.8500 0.0000 1173.9500 0.5200 ;
    END
  END out[216]
  PIN out[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1180.8500 0.0000 1180.9500 0.5200 ;
    END
  END out[215]
  PIN out[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1187.8500 0.0000 1187.9500 0.5200 ;
    END
  END out[214]
  PIN out[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1194.8500 0.0000 1194.9500 0.5200 ;
    END
  END out[213]
  PIN out[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1201.8500 0.0000 1201.9500 0.5200 ;
    END
  END out[212]
  PIN out[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1208.8500 0.0000 1208.9500 0.5200 ;
    END
  END out[211]
  PIN out[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1215.8500 0.0000 1215.9500 0.5200 ;
    END
  END out[210]
  PIN out[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1222.8500 0.0000 1222.9500 0.5200 ;
    END
  END out[209]
  PIN out[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1229.8500 0.0000 1229.9500 0.5200 ;
    END
  END out[208]
  PIN out[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1236.8500 0.0000 1236.9500 0.5200 ;
    END
  END out[207]
  PIN out[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1243.8500 0.0000 1243.9500 0.5200 ;
    END
  END out[206]
  PIN out[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1250.8500 0.0000 1250.9500 0.5200 ;
    END
  END out[205]
  PIN out[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1257.8500 0.0000 1257.9500 0.5200 ;
    END
  END out[204]
  PIN out[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1264.8500 0.0000 1264.9500 0.5200 ;
    END
  END out[203]
  PIN out[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1271.8500 0.0000 1271.9500 0.5200 ;
    END
  END out[202]
  PIN out[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1278.8500 0.0000 1278.9500 0.5200 ;
    END
  END out[201]
  PIN out[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1285.8500 0.0000 1285.9500 0.5200 ;
    END
  END out[200]
  PIN out[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1292.8500 0.0000 1292.9500 0.5200 ;
    END
  END out[199]
  PIN out[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1299.8500 0.0000 1299.9500 0.5200 ;
    END
  END out[198]
  PIN out[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1306.8500 0.0000 1306.9500 0.5200 ;
    END
  END out[197]
  PIN out[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1313.8500 0.0000 1313.9500 0.5200 ;
    END
  END out[196]
  PIN out[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1320.8500 0.0000 1320.9500 0.5200 ;
    END
  END out[195]
  PIN out[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1327.8500 0.0000 1327.9500 0.5200 ;
    END
  END out[194]
  PIN out[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1334.8500 0.0000 1334.9500 0.5200 ;
    END
  END out[193]
  PIN out[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1341.8500 0.0000 1341.9500 0.5200 ;
    END
  END out[192]
  PIN out[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1348.8500 0.0000 1348.9500 0.5200 ;
    END
  END out[191]
  PIN out[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1355.8500 0.0000 1355.9500 0.5200 ;
    END
  END out[190]
  PIN out[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1362.8500 0.0000 1362.9500 0.5200 ;
    END
  END out[189]
  PIN out[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1369.8500 0.0000 1369.9500 0.5200 ;
    END
  END out[188]
  PIN out[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1376.8500 0.0000 1376.9500 0.5200 ;
    END
  END out[187]
  PIN out[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1383.8500 0.0000 1383.9500 0.5200 ;
    END
  END out[186]
  PIN out[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1390.8500 0.0000 1390.9500 0.5200 ;
    END
  END out[185]
  PIN out[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1397.8500 0.0000 1397.9500 0.5200 ;
    END
  END out[184]
  PIN out[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1404.8500 0.0000 1404.9500 0.5200 ;
    END
  END out[183]
  PIN out[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1411.8500 0.0000 1411.9500 0.5200 ;
    END
  END out[182]
  PIN out[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1418.8500 0.0000 1418.9500 0.5200 ;
    END
  END out[181]
  PIN out[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1425.8500 0.0000 1425.9500 0.5200 ;
    END
  END out[180]
  PIN out[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1432.8500 0.0000 1432.9500 0.5200 ;
    END
  END out[179]
  PIN out[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1439.8500 0.0000 1439.9500 0.5200 ;
    END
  END out[178]
  PIN out[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1446.8500 0.0000 1446.9500 0.5200 ;
    END
  END out[177]
  PIN out[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1453.8500 0.0000 1453.9500 0.5200 ;
    END
  END out[176]
  PIN out[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1460.8500 0.0000 1460.9500 0.5200 ;
    END
  END out[175]
  PIN out[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1467.8500 0.0000 1467.9500 0.5200 ;
    END
  END out[174]
  PIN out[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1474.8500 0.0000 1474.9500 0.5200 ;
    END
  END out[173]
  PIN out[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1481.8500 0.0000 1481.9500 0.5200 ;
    END
  END out[172]
  PIN out[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1488.8500 0.0000 1488.9500 0.5200 ;
    END
  END out[171]
  PIN out[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1495.8500 0.0000 1495.9500 0.5200 ;
    END
  END out[170]
  PIN out[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1502.8500 0.0000 1502.9500 0.5200 ;
    END
  END out[169]
  PIN out[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1509.8500 0.0000 1509.9500 0.5200 ;
    END
  END out[168]
  PIN out[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1516.8500 0.0000 1516.9500 0.5200 ;
    END
  END out[167]
  PIN out[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1523.8500 0.0000 1523.9500 0.5200 ;
    END
  END out[166]
  PIN out[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1530.8500 0.0000 1530.9500 0.5200 ;
    END
  END out[165]
  PIN out[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1537.8500 0.0000 1537.9500 0.5200 ;
    END
  END out[164]
  PIN out[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1544.8500 0.0000 1544.9500 0.5200 ;
    END
  END out[163]
  PIN out[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1551.8500 0.0000 1551.9500 0.5200 ;
    END
  END out[162]
  PIN out[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1558.8500 0.0000 1558.9500 0.5200 ;
    END
  END out[161]
  PIN out[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1565.8500 0.0000 1565.9500 0.5200 ;
    END
  END out[160]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 652.0500 0.0000 652.1500 0.5200 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 645.0500 0.0000 645.1500 0.5200 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 638.0500 0.0000 638.1500 0.5200 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 631.0500 0.0000 631.1500 0.5200 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 624.0500 0.0000 624.1500 0.5200 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 617.0500 0.0000 617.1500 0.5200 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 610.0500 0.0000 610.1500 0.5200 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 603.0500 0.0000 603.1500 0.5200 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 596.0500 0.0000 596.1500 0.5200 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 589.0500 0.0000 589.1500 0.5200 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 582.0500 0.0000 582.1500 0.5200 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 575.0500 0.0000 575.1500 0.5200 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 568.0500 0.0000 568.1500 0.5200 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 561.0500 0.0000 561.1500 0.5200 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 554.0500 0.0000 554.1500 0.5200 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 547.0500 0.0000 547.1500 0.5200 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 540.0500 0.0000 540.1500 0.5200 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 533.0500 0.0000 533.1500 0.5200 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 526.0500 0.0000 526.1500 0.5200 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 519.0500 0.0000 519.1500 0.5200 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 512.0500 0.0000 512.1500 0.5200 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 505.0500 0.0000 505.1500 0.5200 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 498.0500 0.0000 498.1500 0.5200 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 491.0500 0.0000 491.1500 0.5200 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 484.0500 0.0000 484.1500 0.5200 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 477.0500 0.0000 477.1500 0.5200 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 470.0500 0.0000 470.1500 0.5200 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 463.0500 0.0000 463.1500 0.5200 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 456.0500 0.0000 456.1500 0.5200 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 449.0500 0.0000 449.1500 0.5200 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 442.0500 0.0000 442.1500 0.5200 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 435.0500 0.0000 435.1500 0.5200 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 428.0500 0.0000 428.1500 0.5200 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 421.0500 0.0000 421.1500 0.5200 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 414.0500 0.0000 414.1500 0.5200 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 407.0500 0.0000 407.1500 0.5200 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 400.0500 0.0000 400.1500 0.5200 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 393.0500 0.0000 393.1500 0.5200 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 386.0500 0.0000 386.1500 0.5200 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 379.0500 0.0000 379.1500 0.5200 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 372.0500 0.0000 372.1500 0.5200 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 365.0500 0.0000 365.1500 0.5200 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 358.0500 0.0000 358.1500 0.5200 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 351.0500 0.0000 351.1500 0.5200 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 344.0500 0.0000 344.1500 0.5200 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 337.0500 0.0000 337.1500 0.5200 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 330.0500 0.0000 330.1500 0.5200 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 323.0500 0.0000 323.1500 0.5200 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 316.0500 0.0000 316.1500 0.5200 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 309.0500 0.0000 309.1500 0.5200 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 302.0500 0.0000 302.1500 0.5200 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 295.0500 0.0000 295.1500 0.5200 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 288.0500 0.0000 288.1500 0.5200 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 281.0500 0.0000 281.1500 0.5200 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 274.0500 0.0000 274.1500 0.5200 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 267.0500 0.0000 267.1500 0.5200 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 260.0500 0.0000 260.1500 0.5200 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 253.0500 0.0000 253.1500 0.5200 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 246.0500 0.0000 246.1500 0.5200 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 239.0500 0.0000 239.1500 0.5200 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 232.0500 0.0000 232.1500 0.5200 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 225.0500 0.0000 225.1500 0.5200 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 218.0500 0.0000 218.1500 0.5200 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 211.0500 0.0000 211.1500 0.5200 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 204.0500 0.0000 204.1500 0.5200 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 197.0500 0.0000 197.1500 0.5200 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 190.0500 0.0000 190.1500 0.5200 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 183.0500 0.0000 183.1500 0.5200 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 176.0500 0.0000 176.1500 0.5200 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 169.0500 0.0000 169.1500 0.5200 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 162.0500 0.0000 162.1500 0.5200 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 155.0500 0.0000 155.1500 0.5200 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 148.0500 0.0000 148.1500 0.5200 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 141.0500 0.0000 141.1500 0.5200 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 134.0500 0.0000 134.1500 0.5200 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 127.0500 0.0000 127.1500 0.5200 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 120.0500 0.0000 120.1500 0.5200 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0500 0.0000 113.1500 0.5200 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 106.0500 0.0000 106.1500 0.5200 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 99.0500 0.0000 99.1500 0.5200 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 648.6500 0.0000 648.7500 0.5200 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 641.6500 0.0000 641.7500 0.5200 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.6500 0.0000 634.7500 0.5200 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 627.6500 0.0000 627.7500 0.5200 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 620.6500 0.0000 620.7500 0.5200 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 613.6500 0.0000 613.7500 0.5200 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 606.6500 0.0000 606.7500 0.5200 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 599.6500 0.0000 599.7500 0.5200 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 592.6500 0.0000 592.7500 0.5200 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 585.6500 0.0000 585.7500 0.5200 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 578.6500 0.0000 578.7500 0.5200 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 571.6500 0.0000 571.7500 0.5200 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 564.6500 0.0000 564.7500 0.5200 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 557.6500 0.0000 557.7500 0.5200 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.6500 0.0000 550.7500 0.5200 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 543.6500 0.0000 543.7500 0.5200 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 536.6500 0.0000 536.7500 0.5200 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 529.6500 0.0000 529.7500 0.5200 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 522.6500 0.0000 522.7500 0.5200 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 515.6500 0.0000 515.7500 0.5200 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 508.6500 0.0000 508.7500 0.5200 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 501.6500 0.0000 501.7500 0.5200 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.6500 0.0000 494.7500 0.5200 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 487.6500 0.0000 487.7500 0.5200 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 480.6500 0.0000 480.7500 0.5200 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 473.6500 0.0000 473.7500 0.5200 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 466.6500 0.0000 466.7500 0.5200 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 459.6500 0.0000 459.7500 0.5200 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 452.6500 0.0000 452.7500 0.5200 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 445.6500 0.0000 445.7500 0.5200 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 438.6500 0.0000 438.7500 0.5200 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 431.6500 0.0000 431.7500 0.5200 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 424.6500 0.0000 424.7500 0.5200 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 417.6500 0.0000 417.7500 0.5200 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 410.6500 0.0000 410.7500 0.5200 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 403.6500 0.0000 403.7500 0.5200 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 396.6500 0.0000 396.7500 0.5200 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 389.6500 0.0000 389.7500 0.5200 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 382.6500 0.0000 382.7500 0.5200 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 375.6500 0.0000 375.7500 0.5200 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 368.6500 0.0000 368.7500 0.5200 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 361.6500 0.0000 361.7500 0.5200 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 354.6500 0.0000 354.7500 0.5200 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 347.6500 0.0000 347.7500 0.5200 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 340.6500 0.0000 340.7500 0.5200 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 333.6500 0.0000 333.7500 0.5200 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 326.6500 0.0000 326.7500 0.5200 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 319.6500 0.0000 319.7500 0.5200 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 312.6500 0.0000 312.7500 0.5200 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 305.6500 0.0000 305.7500 0.5200 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 298.6500 0.0000 298.7500 0.5200 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 291.6500 0.0000 291.7500 0.5200 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 284.6500 0.0000 284.7500 0.5200 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 277.6500 0.0000 277.7500 0.5200 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 270.6500 0.0000 270.7500 0.5200 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 263.6500 0.0000 263.7500 0.5200 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 256.6500 0.0000 256.7500 0.5200 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 249.6500 0.0000 249.7500 0.5200 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 242.6500 0.0000 242.7500 0.5200 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 235.6500 0.0000 235.7500 0.5200 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 228.6500 0.0000 228.7500 0.5200 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 221.6500 0.0000 221.7500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 214.6500 0.0000 214.7500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 207.6500 0.0000 207.7500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 200.6500 0.0000 200.7500 0.5200 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 193.6500 0.0000 193.7500 0.5200 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 186.6500 0.0000 186.7500 0.5200 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 179.6500 0.0000 179.7500 0.5200 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 172.6500 0.0000 172.7500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 165.6500 0.0000 165.7500 0.5200 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 158.6500 0.0000 158.7500 0.5200 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 151.6500 0.0000 151.7500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 144.6500 0.0000 144.7500 0.5200 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 137.6500 0.0000 137.7500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 130.6500 0.0000 130.7500 0.5200 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 123.6500 0.0000 123.7500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 116.6500 0.0000 116.7500 0.5200 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 109.6500 0.0000 109.7500 0.5200 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 102.6500 0.0000 102.7500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 95.6500 0.0000 95.7500 0.5200 ;
    END
  END out[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1761.4000 1760.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 1761.4000 1760.6000 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 1761.4000 1760.6000 ;
    LAYER M4 ;
      RECT 0.0000 0.6200 1761.4000 1760.6000 ;
      RECT 1566.0500 0.0000 1761.4000 0.6200 ;
      RECT 1559.0500 0.0000 1565.7500 0.6200 ;
      RECT 1552.0500 0.0000 1558.7500 0.6200 ;
      RECT 1545.0500 0.0000 1551.7500 0.6200 ;
      RECT 1538.0500 0.0000 1544.7500 0.6200 ;
      RECT 1531.0500 0.0000 1537.7500 0.6200 ;
      RECT 1524.0500 0.0000 1530.7500 0.6200 ;
      RECT 1517.0500 0.0000 1523.7500 0.6200 ;
      RECT 1510.0500 0.0000 1516.7500 0.6200 ;
      RECT 1503.0500 0.0000 1509.7500 0.6200 ;
      RECT 1496.0500 0.0000 1502.7500 0.6200 ;
      RECT 1489.0500 0.0000 1495.7500 0.6200 ;
      RECT 1482.0500 0.0000 1488.7500 0.6200 ;
      RECT 1475.0500 0.0000 1481.7500 0.6200 ;
      RECT 1468.0500 0.0000 1474.7500 0.6200 ;
      RECT 1461.0500 0.0000 1467.7500 0.6200 ;
      RECT 1454.0500 0.0000 1460.7500 0.6200 ;
      RECT 1447.0500 0.0000 1453.7500 0.6200 ;
      RECT 1440.0500 0.0000 1446.7500 0.6200 ;
      RECT 1433.0500 0.0000 1439.7500 0.6200 ;
      RECT 1426.0500 0.0000 1432.7500 0.6200 ;
      RECT 1419.0500 0.0000 1425.7500 0.6200 ;
      RECT 1412.0500 0.0000 1418.7500 0.6200 ;
      RECT 1405.0500 0.0000 1411.7500 0.6200 ;
      RECT 1398.0500 0.0000 1404.7500 0.6200 ;
      RECT 1391.0500 0.0000 1397.7500 0.6200 ;
      RECT 1384.0500 0.0000 1390.7500 0.6200 ;
      RECT 1377.0500 0.0000 1383.7500 0.6200 ;
      RECT 1370.0500 0.0000 1376.7500 0.6200 ;
      RECT 1363.0500 0.0000 1369.7500 0.6200 ;
      RECT 1356.0500 0.0000 1362.7500 0.6200 ;
      RECT 1349.0500 0.0000 1355.7500 0.6200 ;
      RECT 1342.0500 0.0000 1348.7500 0.6200 ;
      RECT 1335.0500 0.0000 1341.7500 0.6200 ;
      RECT 1328.0500 0.0000 1334.7500 0.6200 ;
      RECT 1321.0500 0.0000 1327.7500 0.6200 ;
      RECT 1314.0500 0.0000 1320.7500 0.6200 ;
      RECT 1307.0500 0.0000 1313.7500 0.6200 ;
      RECT 1300.0500 0.0000 1306.7500 0.6200 ;
      RECT 1293.0500 0.0000 1299.7500 0.6200 ;
      RECT 1286.0500 0.0000 1292.7500 0.6200 ;
      RECT 1279.0500 0.0000 1285.7500 0.6200 ;
      RECT 1272.0500 0.0000 1278.7500 0.6200 ;
      RECT 1265.0500 0.0000 1271.7500 0.6200 ;
      RECT 1258.0500 0.0000 1264.7500 0.6200 ;
      RECT 1251.0500 0.0000 1257.7500 0.6200 ;
      RECT 1244.0500 0.0000 1250.7500 0.6200 ;
      RECT 1237.0500 0.0000 1243.7500 0.6200 ;
      RECT 1230.0500 0.0000 1236.7500 0.6200 ;
      RECT 1223.0500 0.0000 1229.7500 0.6200 ;
      RECT 1216.0500 0.0000 1222.7500 0.6200 ;
      RECT 1209.0500 0.0000 1215.7500 0.6200 ;
      RECT 1202.0500 0.0000 1208.7500 0.6200 ;
      RECT 1195.0500 0.0000 1201.7500 0.6200 ;
      RECT 1188.0500 0.0000 1194.7500 0.6200 ;
      RECT 1181.0500 0.0000 1187.7500 0.6200 ;
      RECT 1174.0500 0.0000 1180.7500 0.6200 ;
      RECT 1167.0500 0.0000 1173.7500 0.6200 ;
      RECT 1160.0500 0.0000 1166.7500 0.6200 ;
      RECT 1153.0500 0.0000 1159.7500 0.6200 ;
      RECT 1146.0500 0.0000 1152.7500 0.6200 ;
      RECT 1139.0500 0.0000 1145.7500 0.6200 ;
      RECT 1132.0500 0.0000 1138.7500 0.6200 ;
      RECT 1125.0500 0.0000 1131.7500 0.6200 ;
      RECT 1118.0500 0.0000 1124.7500 0.6200 ;
      RECT 1111.0500 0.0000 1117.7500 0.6200 ;
      RECT 1104.0500 0.0000 1110.7500 0.6200 ;
      RECT 1097.0500 0.0000 1103.7500 0.6200 ;
      RECT 1090.0500 0.0000 1096.7500 0.6200 ;
      RECT 1083.0500 0.0000 1089.7500 0.6200 ;
      RECT 1076.0500 0.0000 1082.7500 0.6200 ;
      RECT 1069.0500 0.0000 1075.7500 0.6200 ;
      RECT 1062.0500 0.0000 1068.7500 0.6200 ;
      RECT 1055.0500 0.0000 1061.7500 0.6200 ;
      RECT 1048.0500 0.0000 1054.7500 0.6200 ;
      RECT 1041.0500 0.0000 1047.7500 0.6200 ;
      RECT 1034.0500 0.0000 1040.7500 0.6200 ;
      RECT 1027.0500 0.0000 1033.7500 0.6200 ;
      RECT 1020.0500 0.0000 1026.7500 0.6200 ;
      RECT 1013.0500 0.0000 1019.7500 0.6200 ;
      RECT 648.8500 0.0000 1012.7500 0.6200 ;
      RECT 641.8500 0.0000 648.5500 0.6200 ;
      RECT 634.8500 0.0000 641.5500 0.6200 ;
      RECT 627.8500 0.0000 634.5500 0.6200 ;
      RECT 620.8500 0.0000 627.5500 0.6200 ;
      RECT 613.8500 0.0000 620.5500 0.6200 ;
      RECT 606.8500 0.0000 613.5500 0.6200 ;
      RECT 599.8500 0.0000 606.5500 0.6200 ;
      RECT 592.8500 0.0000 599.5500 0.6200 ;
      RECT 585.8500 0.0000 592.5500 0.6200 ;
      RECT 578.8500 0.0000 585.5500 0.6200 ;
      RECT 571.8500 0.0000 578.5500 0.6200 ;
      RECT 564.8500 0.0000 571.5500 0.6200 ;
      RECT 557.8500 0.0000 564.5500 0.6200 ;
      RECT 550.8500 0.0000 557.5500 0.6200 ;
      RECT 543.8500 0.0000 550.5500 0.6200 ;
      RECT 536.8500 0.0000 543.5500 0.6200 ;
      RECT 529.8500 0.0000 536.5500 0.6200 ;
      RECT 522.8500 0.0000 529.5500 0.6200 ;
      RECT 515.8500 0.0000 522.5500 0.6200 ;
      RECT 508.8500 0.0000 515.5500 0.6200 ;
      RECT 501.8500 0.0000 508.5500 0.6200 ;
      RECT 494.8500 0.0000 501.5500 0.6200 ;
      RECT 487.8500 0.0000 494.5500 0.6200 ;
      RECT 480.8500 0.0000 487.5500 0.6200 ;
      RECT 473.8500 0.0000 480.5500 0.6200 ;
      RECT 466.8500 0.0000 473.5500 0.6200 ;
      RECT 459.8500 0.0000 466.5500 0.6200 ;
      RECT 452.8500 0.0000 459.5500 0.6200 ;
      RECT 445.8500 0.0000 452.5500 0.6200 ;
      RECT 438.8500 0.0000 445.5500 0.6200 ;
      RECT 431.8500 0.0000 438.5500 0.6200 ;
      RECT 424.8500 0.0000 431.5500 0.6200 ;
      RECT 417.8500 0.0000 424.5500 0.6200 ;
      RECT 410.8500 0.0000 417.5500 0.6200 ;
      RECT 403.8500 0.0000 410.5500 0.6200 ;
      RECT 396.8500 0.0000 403.5500 0.6200 ;
      RECT 389.8500 0.0000 396.5500 0.6200 ;
      RECT 382.8500 0.0000 389.5500 0.6200 ;
      RECT 375.8500 0.0000 382.5500 0.6200 ;
      RECT 368.8500 0.0000 375.5500 0.6200 ;
      RECT 361.8500 0.0000 368.5500 0.6200 ;
      RECT 354.8500 0.0000 361.5500 0.6200 ;
      RECT 347.8500 0.0000 354.5500 0.6200 ;
      RECT 340.8500 0.0000 347.5500 0.6200 ;
      RECT 333.8500 0.0000 340.5500 0.6200 ;
      RECT 326.8500 0.0000 333.5500 0.6200 ;
      RECT 319.8500 0.0000 326.5500 0.6200 ;
      RECT 312.8500 0.0000 319.5500 0.6200 ;
      RECT 305.8500 0.0000 312.5500 0.6200 ;
      RECT 298.8500 0.0000 305.5500 0.6200 ;
      RECT 291.8500 0.0000 298.5500 0.6200 ;
      RECT 284.8500 0.0000 291.5500 0.6200 ;
      RECT 277.8500 0.0000 284.5500 0.6200 ;
      RECT 270.8500 0.0000 277.5500 0.6200 ;
      RECT 263.8500 0.0000 270.5500 0.6200 ;
      RECT 256.8500 0.0000 263.5500 0.6200 ;
      RECT 249.8500 0.0000 256.5500 0.6200 ;
      RECT 242.8500 0.0000 249.5500 0.6200 ;
      RECT 235.8500 0.0000 242.5500 0.6200 ;
      RECT 228.8500 0.0000 235.5500 0.6200 ;
      RECT 221.8500 0.0000 228.5500 0.6200 ;
      RECT 214.8500 0.0000 221.5500 0.6200 ;
      RECT 207.8500 0.0000 214.5500 0.6200 ;
      RECT 200.8500 0.0000 207.5500 0.6200 ;
      RECT 193.8500 0.0000 200.5500 0.6200 ;
      RECT 186.8500 0.0000 193.5500 0.6200 ;
      RECT 179.8500 0.0000 186.5500 0.6200 ;
      RECT 172.8500 0.0000 179.5500 0.6200 ;
      RECT 165.8500 0.0000 172.5500 0.6200 ;
      RECT 158.8500 0.0000 165.5500 0.6200 ;
      RECT 151.8500 0.0000 158.5500 0.6200 ;
      RECT 144.8500 0.0000 151.5500 0.6200 ;
      RECT 137.8500 0.0000 144.5500 0.6200 ;
      RECT 130.8500 0.0000 137.5500 0.6200 ;
      RECT 123.8500 0.0000 130.5500 0.6200 ;
      RECT 116.8500 0.0000 123.5500 0.6200 ;
      RECT 109.8500 0.0000 116.5500 0.6200 ;
      RECT 102.8500 0.0000 109.5500 0.6200 ;
      RECT 95.8500 0.0000 102.5500 0.6200 ;
      RECT 0.0000 0.0000 95.5500 0.6200 ;
    LAYER M5 ;
      RECT 0.0000 669.1500 1761.4000 1760.6000 ;
      RECT 0.6200 668.8500 1760.7800 669.1500 ;
      RECT 0.0000 665.1500 1761.4000 668.8500 ;
      RECT 0.6200 664.8500 1760.7800 665.1500 ;
      RECT 0.0000 661.1500 1761.4000 664.8500 ;
      RECT 0.6200 660.8500 1760.7800 661.1500 ;
      RECT 0.0000 657.1500 1761.4000 660.8500 ;
      RECT 0.6200 656.8500 1760.7800 657.1500 ;
      RECT 0.0000 653.1500 1761.4000 656.8500 ;
      RECT 0.6200 652.8500 1760.7800 653.1500 ;
      RECT 0.0000 649.1500 1761.4000 652.8500 ;
      RECT 0.6200 648.8500 1760.7800 649.1500 ;
      RECT 0.0000 645.1500 1761.4000 648.8500 ;
      RECT 0.6200 644.8500 1760.7800 645.1500 ;
      RECT 0.0000 641.1500 1761.4000 644.8500 ;
      RECT 0.6200 640.8500 1760.7800 641.1500 ;
      RECT 0.0000 637.1500 1761.4000 640.8500 ;
      RECT 0.6200 636.8500 1760.7800 637.1500 ;
      RECT 0.0000 633.1500 1761.4000 636.8500 ;
      RECT 0.6200 632.8500 1760.7800 633.1500 ;
      RECT 0.0000 629.1500 1761.4000 632.8500 ;
      RECT 0.6200 628.8500 1760.7800 629.1500 ;
      RECT 0.0000 625.1500 1761.4000 628.8500 ;
      RECT 0.6200 624.8500 1760.7800 625.1500 ;
      RECT 0.0000 621.1500 1761.4000 624.8500 ;
      RECT 0.6200 620.8500 1760.7800 621.1500 ;
      RECT 0.0000 617.1500 1761.4000 620.8500 ;
      RECT 0.6200 616.8500 1760.7800 617.1500 ;
      RECT 0.0000 613.1500 1761.4000 616.8500 ;
      RECT 0.6200 612.8500 1760.7800 613.1500 ;
      RECT 0.0000 609.1500 1761.4000 612.8500 ;
      RECT 0.6200 608.8500 1760.7800 609.1500 ;
      RECT 0.0000 605.1500 1761.4000 608.8500 ;
      RECT 0.6200 604.8500 1760.7800 605.1500 ;
      RECT 0.0000 601.1500 1761.4000 604.8500 ;
      RECT 0.6200 600.8500 1760.7800 601.1500 ;
      RECT 0.0000 597.1500 1761.4000 600.8500 ;
      RECT 0.6200 596.8500 1760.7800 597.1500 ;
      RECT 0.0000 593.1500 1761.4000 596.8500 ;
      RECT 0.6200 592.8500 1760.7800 593.1500 ;
      RECT 0.0000 589.1500 1761.4000 592.8500 ;
      RECT 0.6200 588.8500 1760.7800 589.1500 ;
      RECT 0.0000 585.1500 1761.4000 588.8500 ;
      RECT 0.6200 584.8500 1760.7800 585.1500 ;
      RECT 0.0000 581.1500 1761.4000 584.8500 ;
      RECT 0.6200 580.8500 1760.7800 581.1500 ;
      RECT 0.0000 577.1500 1761.4000 580.8500 ;
      RECT 0.6200 576.8500 1760.7800 577.1500 ;
      RECT 0.0000 573.1500 1761.4000 576.8500 ;
      RECT 0.6200 572.8500 1760.7800 573.1500 ;
      RECT 0.0000 569.1500 1761.4000 572.8500 ;
      RECT 0.6200 568.8500 1760.7800 569.1500 ;
      RECT 0.0000 565.1500 1761.4000 568.8500 ;
      RECT 0.6200 564.8500 1760.7800 565.1500 ;
      RECT 0.0000 561.1500 1761.4000 564.8500 ;
      RECT 0.6200 560.8500 1760.7800 561.1500 ;
      RECT 0.0000 557.1500 1761.4000 560.8500 ;
      RECT 0.6200 556.8500 1760.7800 557.1500 ;
      RECT 0.0000 553.1500 1761.4000 556.8500 ;
      RECT 0.6200 552.8500 1760.7800 553.1500 ;
      RECT 0.0000 549.1500 1761.4000 552.8500 ;
      RECT 0.6200 548.8500 1760.7800 549.1500 ;
      RECT 0.0000 545.1500 1761.4000 548.8500 ;
      RECT 0.6200 544.8500 1760.7800 545.1500 ;
      RECT 0.0000 541.1500 1761.4000 544.8500 ;
      RECT 0.6200 540.8500 1760.7800 541.1500 ;
      RECT 0.0000 537.1500 1761.4000 540.8500 ;
      RECT 0.6200 536.8500 1760.7800 537.1500 ;
      RECT 0.0000 533.1500 1761.4000 536.8500 ;
      RECT 0.6200 532.8500 1760.7800 533.1500 ;
      RECT 0.0000 529.1500 1761.4000 532.8500 ;
      RECT 0.6200 528.8500 1760.7800 529.1500 ;
      RECT 0.0000 525.1500 1761.4000 528.8500 ;
      RECT 0.6200 524.8500 1760.7800 525.1500 ;
      RECT 0.0000 521.1500 1761.4000 524.8500 ;
      RECT 0.6200 520.8500 1760.7800 521.1500 ;
      RECT 0.0000 517.1500 1761.4000 520.8500 ;
      RECT 0.6200 516.8500 1760.7800 517.1500 ;
      RECT 0.0000 513.1500 1761.4000 516.8500 ;
      RECT 0.6200 512.8500 1760.7800 513.1500 ;
      RECT 0.0000 509.1500 1761.4000 512.8500 ;
      RECT 0.6200 508.8500 1760.7800 509.1500 ;
      RECT 0.0000 505.1500 1761.4000 508.8500 ;
      RECT 0.6200 504.8500 1760.7800 505.1500 ;
      RECT 0.0000 501.1500 1761.4000 504.8500 ;
      RECT 0.6200 500.8500 1760.7800 501.1500 ;
      RECT 0.0000 497.1500 1761.4000 500.8500 ;
      RECT 0.6200 496.8500 1760.7800 497.1500 ;
      RECT 0.0000 493.1500 1761.4000 496.8500 ;
      RECT 0.6200 492.8500 1760.7800 493.1500 ;
      RECT 0.0000 489.1500 1761.4000 492.8500 ;
      RECT 0.6200 488.8500 1760.7800 489.1500 ;
      RECT 0.0000 485.1500 1761.4000 488.8500 ;
      RECT 0.6200 484.8500 1760.7800 485.1500 ;
      RECT 0.0000 481.1500 1761.4000 484.8500 ;
      RECT 0.6200 480.8500 1760.7800 481.1500 ;
      RECT 0.0000 477.1500 1761.4000 480.8500 ;
      RECT 0.6200 476.8500 1760.7800 477.1500 ;
      RECT 0.0000 473.1500 1761.4000 476.8500 ;
      RECT 0.6200 472.8500 1760.7800 473.1500 ;
      RECT 0.0000 469.1500 1761.4000 472.8500 ;
      RECT 0.6200 468.8500 1760.7800 469.1500 ;
      RECT 0.0000 465.1500 1761.4000 468.8500 ;
      RECT 0.6200 464.8500 1760.7800 465.1500 ;
      RECT 0.0000 461.1500 1761.4000 464.8500 ;
      RECT 0.6200 460.8500 1760.7800 461.1500 ;
      RECT 0.0000 457.1500 1761.4000 460.8500 ;
      RECT 0.6200 456.8500 1760.7800 457.1500 ;
      RECT 0.0000 453.1500 1761.4000 456.8500 ;
      RECT 0.6200 452.8500 1760.7800 453.1500 ;
      RECT 0.0000 449.1500 1761.4000 452.8500 ;
      RECT 0.6200 448.8500 1760.7800 449.1500 ;
      RECT 0.0000 445.1500 1761.4000 448.8500 ;
      RECT 0.6200 444.8500 1760.7800 445.1500 ;
      RECT 0.0000 441.1500 1761.4000 444.8500 ;
      RECT 0.6200 440.8500 1760.7800 441.1500 ;
      RECT 0.0000 437.1500 1761.4000 440.8500 ;
      RECT 0.6200 436.8500 1760.7800 437.1500 ;
      RECT 0.0000 433.1500 1761.4000 436.8500 ;
      RECT 0.6200 432.8500 1760.7800 433.1500 ;
      RECT 0.0000 429.1500 1761.4000 432.8500 ;
      RECT 0.6200 428.8500 1760.7800 429.1500 ;
      RECT 0.0000 425.1500 1761.4000 428.8500 ;
      RECT 0.6200 424.8500 1760.7800 425.1500 ;
      RECT 0.0000 421.1500 1761.4000 424.8500 ;
      RECT 0.6200 420.8500 1760.7800 421.1500 ;
      RECT 0.0000 417.1500 1761.4000 420.8500 ;
      RECT 0.6200 416.8500 1760.7800 417.1500 ;
      RECT 0.0000 413.1500 1761.4000 416.8500 ;
      RECT 0.6200 412.8500 1760.7800 413.1500 ;
      RECT 0.0000 409.1500 1761.4000 412.8500 ;
      RECT 0.6200 408.8500 1760.7800 409.1500 ;
      RECT 0.0000 405.1500 1761.4000 408.8500 ;
      RECT 0.6200 404.8500 1760.7800 405.1500 ;
      RECT 0.0000 401.1500 1761.4000 404.8500 ;
      RECT 0.6200 400.8500 1760.7800 401.1500 ;
      RECT 0.0000 397.1500 1761.4000 400.8500 ;
      RECT 0.6200 396.8500 1760.7800 397.1500 ;
      RECT 0.0000 393.1500 1761.4000 396.8500 ;
      RECT 0.6200 392.8500 1760.7800 393.1500 ;
      RECT 0.0000 389.1500 1761.4000 392.8500 ;
      RECT 0.6200 388.8500 1760.7800 389.1500 ;
      RECT 0.0000 385.1500 1761.4000 388.8500 ;
      RECT 0.6200 384.8500 1760.7800 385.1500 ;
      RECT 0.0000 381.1500 1761.4000 384.8500 ;
      RECT 0.6200 380.8500 1760.7800 381.1500 ;
      RECT 0.0000 377.1500 1761.4000 380.8500 ;
      RECT 0.6200 376.8500 1760.7800 377.1500 ;
      RECT 0.0000 373.1500 1761.4000 376.8500 ;
      RECT 0.6200 372.8500 1760.7800 373.1500 ;
      RECT 0.0000 369.1500 1761.4000 372.8500 ;
      RECT 0.6200 368.8500 1760.7800 369.1500 ;
      RECT 0.0000 365.1500 1761.4000 368.8500 ;
      RECT 0.6200 364.8500 1760.7800 365.1500 ;
      RECT 0.0000 361.1500 1761.4000 364.8500 ;
      RECT 0.6200 360.8500 1760.7800 361.1500 ;
      RECT 0.0000 357.1500 1761.4000 360.8500 ;
      RECT 0.6200 356.8500 1760.7800 357.1500 ;
      RECT 0.0000 353.1500 1761.4000 356.8500 ;
      RECT 0.6200 352.8500 1760.7800 353.1500 ;
      RECT 0.0000 349.1500 1761.4000 352.8500 ;
      RECT 0.6200 348.8500 1760.7800 349.1500 ;
      RECT 0.0000 345.1500 1761.4000 348.8500 ;
      RECT 0.6200 344.8500 1760.7800 345.1500 ;
      RECT 0.0000 341.1500 1761.4000 344.8500 ;
      RECT 0.6200 340.8500 1760.7800 341.1500 ;
      RECT 0.0000 337.1500 1761.4000 340.8500 ;
      RECT 0.6200 336.8500 1760.7800 337.1500 ;
      RECT 0.0000 333.1500 1761.4000 336.8500 ;
      RECT 0.6200 332.8500 1760.7800 333.1500 ;
      RECT 0.0000 329.1500 1761.4000 332.8500 ;
      RECT 0.6200 328.8500 1760.7800 329.1500 ;
      RECT 0.0000 325.1500 1761.4000 328.8500 ;
      RECT 0.6200 324.8500 1760.7800 325.1500 ;
      RECT 0.0000 0.0000 1761.4000 324.8500 ;
    LAYER M6 ;
      RECT 0.0000 0.6200 1761.4000 1760.6000 ;
      RECT 1562.6500 0.0000 1761.4000 0.6200 ;
      RECT 1555.6500 0.0000 1562.3500 0.6200 ;
      RECT 1548.6500 0.0000 1555.3500 0.6200 ;
      RECT 1541.6500 0.0000 1548.3500 0.6200 ;
      RECT 1534.6500 0.0000 1541.3500 0.6200 ;
      RECT 1527.6500 0.0000 1534.3500 0.6200 ;
      RECT 1520.6500 0.0000 1527.3500 0.6200 ;
      RECT 1513.6500 0.0000 1520.3500 0.6200 ;
      RECT 1506.6500 0.0000 1513.3500 0.6200 ;
      RECT 1499.6500 0.0000 1506.3500 0.6200 ;
      RECT 1492.6500 0.0000 1499.3500 0.6200 ;
      RECT 1485.6500 0.0000 1492.3500 0.6200 ;
      RECT 1478.6500 0.0000 1485.3500 0.6200 ;
      RECT 1471.6500 0.0000 1478.3500 0.6200 ;
      RECT 1464.6500 0.0000 1471.3500 0.6200 ;
      RECT 1457.6500 0.0000 1464.3500 0.6200 ;
      RECT 1450.6500 0.0000 1457.3500 0.6200 ;
      RECT 1443.6500 0.0000 1450.3500 0.6200 ;
      RECT 1436.6500 0.0000 1443.3500 0.6200 ;
      RECT 1429.6500 0.0000 1436.3500 0.6200 ;
      RECT 1422.6500 0.0000 1429.3500 0.6200 ;
      RECT 1415.6500 0.0000 1422.3500 0.6200 ;
      RECT 1408.6500 0.0000 1415.3500 0.6200 ;
      RECT 1401.6500 0.0000 1408.3500 0.6200 ;
      RECT 1394.6500 0.0000 1401.3500 0.6200 ;
      RECT 1387.6500 0.0000 1394.3500 0.6200 ;
      RECT 1380.6500 0.0000 1387.3500 0.6200 ;
      RECT 1373.6500 0.0000 1380.3500 0.6200 ;
      RECT 1366.6500 0.0000 1373.3500 0.6200 ;
      RECT 1359.6500 0.0000 1366.3500 0.6200 ;
      RECT 1352.6500 0.0000 1359.3500 0.6200 ;
      RECT 1345.6500 0.0000 1352.3500 0.6200 ;
      RECT 1338.6500 0.0000 1345.3500 0.6200 ;
      RECT 1331.6500 0.0000 1338.3500 0.6200 ;
      RECT 1324.6500 0.0000 1331.3500 0.6200 ;
      RECT 1317.6500 0.0000 1324.3500 0.6200 ;
      RECT 1310.6500 0.0000 1317.3500 0.6200 ;
      RECT 1303.6500 0.0000 1310.3500 0.6200 ;
      RECT 1296.6500 0.0000 1303.3500 0.6200 ;
      RECT 1289.6500 0.0000 1296.3500 0.6200 ;
      RECT 1282.6500 0.0000 1289.3500 0.6200 ;
      RECT 1275.6500 0.0000 1282.3500 0.6200 ;
      RECT 1268.6500 0.0000 1275.3500 0.6200 ;
      RECT 1261.6500 0.0000 1268.3500 0.6200 ;
      RECT 1254.6500 0.0000 1261.3500 0.6200 ;
      RECT 1247.6500 0.0000 1254.3500 0.6200 ;
      RECT 1240.6500 0.0000 1247.3500 0.6200 ;
      RECT 1233.6500 0.0000 1240.3500 0.6200 ;
      RECT 1226.6500 0.0000 1233.3500 0.6200 ;
      RECT 1219.6500 0.0000 1226.3500 0.6200 ;
      RECT 1212.6500 0.0000 1219.3500 0.6200 ;
      RECT 1205.6500 0.0000 1212.3500 0.6200 ;
      RECT 1198.6500 0.0000 1205.3500 0.6200 ;
      RECT 1191.6500 0.0000 1198.3500 0.6200 ;
      RECT 1184.6500 0.0000 1191.3500 0.6200 ;
      RECT 1177.6500 0.0000 1184.3500 0.6200 ;
      RECT 1170.6500 0.0000 1177.3500 0.6200 ;
      RECT 1163.6500 0.0000 1170.3500 0.6200 ;
      RECT 1156.6500 0.0000 1163.3500 0.6200 ;
      RECT 1149.6500 0.0000 1156.3500 0.6200 ;
      RECT 1142.6500 0.0000 1149.3500 0.6200 ;
      RECT 1135.6500 0.0000 1142.3500 0.6200 ;
      RECT 1128.6500 0.0000 1135.3500 0.6200 ;
      RECT 1121.6500 0.0000 1128.3500 0.6200 ;
      RECT 1114.6500 0.0000 1121.3500 0.6200 ;
      RECT 1107.6500 0.0000 1114.3500 0.6200 ;
      RECT 1100.6500 0.0000 1107.3500 0.6200 ;
      RECT 1093.6500 0.0000 1100.3500 0.6200 ;
      RECT 1086.6500 0.0000 1093.3500 0.6200 ;
      RECT 1079.6500 0.0000 1086.3500 0.6200 ;
      RECT 1072.6500 0.0000 1079.3500 0.6200 ;
      RECT 1065.6500 0.0000 1072.3500 0.6200 ;
      RECT 1058.6500 0.0000 1065.3500 0.6200 ;
      RECT 1051.6500 0.0000 1058.3500 0.6200 ;
      RECT 1044.6500 0.0000 1051.3500 0.6200 ;
      RECT 1037.6500 0.0000 1044.3500 0.6200 ;
      RECT 1030.6500 0.0000 1037.3500 0.6200 ;
      RECT 1023.6500 0.0000 1030.3500 0.6200 ;
      RECT 1016.6500 0.0000 1023.3500 0.6200 ;
      RECT 1009.6500 0.0000 1016.3500 0.6200 ;
      RECT 881.0500 0.0000 1009.3500 0.6200 ;
      RECT 652.2500 0.0000 880.7500 0.6200 ;
      RECT 645.2500 0.0000 651.9500 0.6200 ;
      RECT 638.2500 0.0000 644.9500 0.6200 ;
      RECT 631.2500 0.0000 637.9500 0.6200 ;
      RECT 624.2500 0.0000 630.9500 0.6200 ;
      RECT 617.2500 0.0000 623.9500 0.6200 ;
      RECT 610.2500 0.0000 616.9500 0.6200 ;
      RECT 603.2500 0.0000 609.9500 0.6200 ;
      RECT 596.2500 0.0000 602.9500 0.6200 ;
      RECT 589.2500 0.0000 595.9500 0.6200 ;
      RECT 582.2500 0.0000 588.9500 0.6200 ;
      RECT 575.2500 0.0000 581.9500 0.6200 ;
      RECT 568.2500 0.0000 574.9500 0.6200 ;
      RECT 561.2500 0.0000 567.9500 0.6200 ;
      RECT 554.2500 0.0000 560.9500 0.6200 ;
      RECT 547.2500 0.0000 553.9500 0.6200 ;
      RECT 540.2500 0.0000 546.9500 0.6200 ;
      RECT 533.2500 0.0000 539.9500 0.6200 ;
      RECT 526.2500 0.0000 532.9500 0.6200 ;
      RECT 519.2500 0.0000 525.9500 0.6200 ;
      RECT 512.2500 0.0000 518.9500 0.6200 ;
      RECT 505.2500 0.0000 511.9500 0.6200 ;
      RECT 498.2500 0.0000 504.9500 0.6200 ;
      RECT 491.2500 0.0000 497.9500 0.6200 ;
      RECT 484.2500 0.0000 490.9500 0.6200 ;
      RECT 477.2500 0.0000 483.9500 0.6200 ;
      RECT 470.2500 0.0000 476.9500 0.6200 ;
      RECT 463.2500 0.0000 469.9500 0.6200 ;
      RECT 456.2500 0.0000 462.9500 0.6200 ;
      RECT 449.2500 0.0000 455.9500 0.6200 ;
      RECT 442.2500 0.0000 448.9500 0.6200 ;
      RECT 435.2500 0.0000 441.9500 0.6200 ;
      RECT 428.2500 0.0000 434.9500 0.6200 ;
      RECT 421.2500 0.0000 427.9500 0.6200 ;
      RECT 414.2500 0.0000 420.9500 0.6200 ;
      RECT 407.2500 0.0000 413.9500 0.6200 ;
      RECT 400.2500 0.0000 406.9500 0.6200 ;
      RECT 393.2500 0.0000 399.9500 0.6200 ;
      RECT 386.2500 0.0000 392.9500 0.6200 ;
      RECT 379.2500 0.0000 385.9500 0.6200 ;
      RECT 372.2500 0.0000 378.9500 0.6200 ;
      RECT 365.2500 0.0000 371.9500 0.6200 ;
      RECT 358.2500 0.0000 364.9500 0.6200 ;
      RECT 351.2500 0.0000 357.9500 0.6200 ;
      RECT 344.2500 0.0000 350.9500 0.6200 ;
      RECT 337.2500 0.0000 343.9500 0.6200 ;
      RECT 330.2500 0.0000 336.9500 0.6200 ;
      RECT 323.2500 0.0000 329.9500 0.6200 ;
      RECT 316.2500 0.0000 322.9500 0.6200 ;
      RECT 309.2500 0.0000 315.9500 0.6200 ;
      RECT 302.2500 0.0000 308.9500 0.6200 ;
      RECT 295.2500 0.0000 301.9500 0.6200 ;
      RECT 288.2500 0.0000 294.9500 0.6200 ;
      RECT 281.2500 0.0000 287.9500 0.6200 ;
      RECT 274.2500 0.0000 280.9500 0.6200 ;
      RECT 267.2500 0.0000 273.9500 0.6200 ;
      RECT 260.2500 0.0000 266.9500 0.6200 ;
      RECT 253.2500 0.0000 259.9500 0.6200 ;
      RECT 246.2500 0.0000 252.9500 0.6200 ;
      RECT 239.2500 0.0000 245.9500 0.6200 ;
      RECT 232.2500 0.0000 238.9500 0.6200 ;
      RECT 225.2500 0.0000 231.9500 0.6200 ;
      RECT 218.2500 0.0000 224.9500 0.6200 ;
      RECT 211.2500 0.0000 217.9500 0.6200 ;
      RECT 204.2500 0.0000 210.9500 0.6200 ;
      RECT 197.2500 0.0000 203.9500 0.6200 ;
      RECT 190.2500 0.0000 196.9500 0.6200 ;
      RECT 183.2500 0.0000 189.9500 0.6200 ;
      RECT 176.2500 0.0000 182.9500 0.6200 ;
      RECT 169.2500 0.0000 175.9500 0.6200 ;
      RECT 162.2500 0.0000 168.9500 0.6200 ;
      RECT 155.2500 0.0000 161.9500 0.6200 ;
      RECT 148.2500 0.0000 154.9500 0.6200 ;
      RECT 141.2500 0.0000 147.9500 0.6200 ;
      RECT 134.2500 0.0000 140.9500 0.6200 ;
      RECT 127.2500 0.0000 133.9500 0.6200 ;
      RECT 120.2500 0.0000 126.9500 0.6200 ;
      RECT 113.2500 0.0000 119.9500 0.6200 ;
      RECT 106.2500 0.0000 112.9500 0.6200 ;
      RECT 99.2500 0.0000 105.9500 0.6200 ;
      RECT 0.0000 0.0000 98.9500 0.6200 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 1761.4000 1760.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 1761.4000 1760.6000 ;
  END
END fullchip

END LIBRARY
