/home/linux/ieng6/ee260bwi25/mak025/ECE260B_Project/single_core/pnr/core/subckt/sram_w8_64b.lef