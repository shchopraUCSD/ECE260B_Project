/home/linux/ieng6/ee260bwi25/sparanjpay/ECE260B_Project/dual_core/pnr/dual_core/subckt/core.lef