##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Wed Mar 19 18:39:00 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w8_64b
  CLASS BLOCK ;
  SIZE 116.4000 BY 115.6000 ;
  FOREIGN sram_w8_64b 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.9500 0.6000 46.0500 ;
    END
  END CLK
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.4500 0.0000 89.5500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4500 0.0000 88.5500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.4500 0.0000 87.5500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.4500 0.0000 86.5500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4500 0.0000 85.5500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.4500 0.0000 84.5500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.4500 0.0000 83.5500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.4500 0.0000 82.5500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.4500 0.0000 81.5500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.4500 0.0000 80.5500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.4500 0.0000 79.5500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.4500 0.0000 78.5500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.4500 0.0000 77.5500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4500 0.0000 76.5500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.4500 0.0000 75.5500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.4500 0.0000 74.5500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.4500 0.0000 73.5500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.4500 0.0000 72.5500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.4500 0.0000 71.5500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.4500 0.0000 70.5500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.4500 0.0000 69.5500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.4500 0.0000 68.5500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.4500 0.0000 67.5500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.4500 0.0000 66.5500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.4500 0.0000 65.5500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4500 0.0000 64.5500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.4500 0.0000 63.5500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.4500 0.0000 62.5500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4500 0.0000 61.5500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.4500 0.0000 60.5500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.4500 0.0000 59.5500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.4500 0.0000 58.5500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.4500 0.0000 57.5500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.4500 0.0000 56.5500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.4500 0.0000 55.5500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.4500 0.0000 54.5500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.4500 0.0000 53.5500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4500 0.0000 52.5500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.4500 0.0000 51.5500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.4500 0.0000 50.5500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.4500 0.0000 49.5500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.4500 0.0000 48.5500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.4500 0.0000 47.5500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4500 0.0000 46.5500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.4500 0.0000 45.5500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.4500 0.0000 44.5500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4500 0.0000 43.5500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.4500 0.0000 42.5500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.4500 0.0000 41.5500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4500 0.0000 40.5500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.4500 0.0000 39.5500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.4500 0.0000 38.5500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4500 0.0000 37.5500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.4500 0.0000 36.5500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.4500 0.0000 35.5500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.4500 0.0000 34.5500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.4500 0.0000 33.5500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4500 0.0000 32.5500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.4500 0.0000 31.5500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.4500 0.0000 30.5500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.4500 0.0000 29.5500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4500 0.0000 28.5500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.4500 0.0000 27.5500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.4500 0.0000 26.5500 0.6000 ;
    END
  END D[0]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.4500 115.0000 89.5500 115.6000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.4500 115.0000 88.5500 115.6000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.4500 115.0000 87.5500 115.6000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.4500 115.0000 86.5500 115.6000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4500 115.0000 85.5500 115.6000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.4500 115.0000 84.5500 115.6000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.4500 115.0000 83.5500 115.6000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.4500 115.0000 82.5500 115.6000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.4500 115.0000 81.5500 115.6000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.4500 115.0000 80.5500 115.6000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.4500 115.0000 79.5500 115.6000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.4500 115.0000 78.5500 115.6000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.4500 115.0000 77.5500 115.6000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.4500 115.0000 76.5500 115.6000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.4500 115.0000 75.5500 115.6000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.4500 115.0000 74.5500 115.6000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.4500 115.0000 73.5500 115.6000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.4500 115.0000 72.5500 115.6000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.4500 115.0000 71.5500 115.6000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.4500 115.0000 70.5500 115.6000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.4500 115.0000 69.5500 115.6000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.4500 115.0000 68.5500 115.6000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.4500 115.0000 67.5500 115.6000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.4500 115.0000 66.5500 115.6000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.4500 115.0000 65.5500 115.6000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.4500 115.0000 64.5500 115.6000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.4500 115.0000 63.5500 115.6000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.4500 115.0000 62.5500 115.6000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4500 115.0000 61.5500 115.6000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.4500 115.0000 60.5500 115.6000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.4500 115.0000 59.5500 115.6000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.4500 115.0000 58.5500 115.6000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.4500 115.0000 57.5500 115.6000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.4500 115.0000 56.5500 115.6000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.4500 115.0000 55.5500 115.6000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.4500 115.0000 54.5500 115.6000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.4500 115.0000 53.5500 115.6000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.4500 115.0000 52.5500 115.6000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.4500 115.0000 51.5500 115.6000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.4500 115.0000 50.5500 115.6000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.4500 115.0000 49.5500 115.6000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.4500 115.0000 48.5500 115.6000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.4500 115.0000 47.5500 115.6000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.4500 115.0000 46.5500 115.6000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.4500 115.0000 45.5500 115.6000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.4500 115.0000 44.5500 115.6000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.4500 115.0000 43.5500 115.6000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.4500 115.0000 42.5500 115.6000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.4500 115.0000 41.5500 115.6000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.4500 115.0000 40.5500 115.6000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.4500 115.0000 39.5500 115.6000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.4500 115.0000 38.5500 115.6000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4500 115.0000 37.5500 115.6000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.4500 115.0000 36.5500 115.6000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.4500 115.0000 35.5500 115.6000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.4500 115.0000 34.5500 115.6000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.4500 115.0000 33.5500 115.6000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.4500 115.0000 32.5500 115.6000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.4500 115.0000 31.5500 115.6000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.4500 115.0000 30.5500 115.6000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.4500 115.0000 29.5500 115.6000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.4500 115.0000 28.5500 115.6000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.4500 115.0000 27.5500 115.6000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.4500 115.0000 26.5500 115.6000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.9500 0.6000 54.0500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.9500 0.6000 50.0500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.9500 0.6000 58.0500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.9500 0.6000 62.0500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.9500 0.6000 66.0500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.9500 0.6000 70.0500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 12.0000 2.0000 14.0000 113.6000 ;
        RECT 28.2200 2.0000 30.2200 113.6000 ;
        RECT 44.4400 2.0000 46.4400 113.6000 ;
        RECT 76.8800 2.0000 78.8800 113.6000 ;
        RECT 60.6600 2.0000 62.6600 113.6000 ;
        RECT 109.3200 2.0000 111.3200 113.6000 ;
        RECT 93.1000 2.0000 95.1000 113.6000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 5.0000 2.0000 7.0000 113.6000 ;
        RECT 21.2200 2.0000 23.2200 113.6000 ;
        RECT 37.4400 2.0000 39.4400 113.6000 ;
        RECT 53.6600 2.0000 55.6600 113.6000 ;
        RECT 86.1000 2.0000 88.1000 113.6000 ;
        RECT 69.8800 2.0000 71.8800 113.6000 ;
        RECT 102.3200 2.0000 104.3200 113.6000 ;
        RECT 5.0000 1.8350 7.0000 2.1650 ;
        RECT 21.2200 1.8350 23.2200 2.1650 ;
        RECT 37.4400 1.8350 39.4400 2.1650 ;
        RECT 53.6600 1.8350 55.6600 2.1650 ;
        RECT 86.1000 1.8350 88.1000 2.1650 ;
        RECT 69.8800 1.8350 71.8800 2.1650 ;
        RECT 102.3200 1.8350 104.3200 2.1650 ;
        RECT 5.0000 113.4350 7.0000 113.7650 ;
        RECT 21.2200 113.4350 23.2200 113.7650 ;
        RECT 37.4400 113.4350 39.4400 113.7650 ;
        RECT 53.6600 113.4350 55.6600 113.7650 ;
        RECT 86.1000 113.4350 88.1000 113.7650 ;
        RECT 69.8800 113.4350 71.8800 113.7650 ;
        RECT 102.3200 113.4350 104.3200 113.7650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 116.4000 115.6000 ;
    LAYER M2 ;
      RECT 89.6500 114.9000 116.4000 115.6000 ;
      RECT 88.6500 114.9000 89.3500 115.6000 ;
      RECT 87.6500 114.9000 88.3500 115.6000 ;
      RECT 86.6500 114.9000 87.3500 115.6000 ;
      RECT 85.6500 114.9000 86.3500 115.6000 ;
      RECT 84.6500 114.9000 85.3500 115.6000 ;
      RECT 83.6500 114.9000 84.3500 115.6000 ;
      RECT 82.6500 114.9000 83.3500 115.6000 ;
      RECT 81.6500 114.9000 82.3500 115.6000 ;
      RECT 80.6500 114.9000 81.3500 115.6000 ;
      RECT 79.6500 114.9000 80.3500 115.6000 ;
      RECT 78.6500 114.9000 79.3500 115.6000 ;
      RECT 77.6500 114.9000 78.3500 115.6000 ;
      RECT 76.6500 114.9000 77.3500 115.6000 ;
      RECT 75.6500 114.9000 76.3500 115.6000 ;
      RECT 74.6500 114.9000 75.3500 115.6000 ;
      RECT 73.6500 114.9000 74.3500 115.6000 ;
      RECT 72.6500 114.9000 73.3500 115.6000 ;
      RECT 71.6500 114.9000 72.3500 115.6000 ;
      RECT 70.6500 114.9000 71.3500 115.6000 ;
      RECT 69.6500 114.9000 70.3500 115.6000 ;
      RECT 68.6500 114.9000 69.3500 115.6000 ;
      RECT 67.6500 114.9000 68.3500 115.6000 ;
      RECT 66.6500 114.9000 67.3500 115.6000 ;
      RECT 65.6500 114.9000 66.3500 115.6000 ;
      RECT 64.6500 114.9000 65.3500 115.6000 ;
      RECT 63.6500 114.9000 64.3500 115.6000 ;
      RECT 62.6500 114.9000 63.3500 115.6000 ;
      RECT 61.6500 114.9000 62.3500 115.6000 ;
      RECT 60.6500 114.9000 61.3500 115.6000 ;
      RECT 59.6500 114.9000 60.3500 115.6000 ;
      RECT 58.6500 114.9000 59.3500 115.6000 ;
      RECT 57.6500 114.9000 58.3500 115.6000 ;
      RECT 56.6500 114.9000 57.3500 115.6000 ;
      RECT 55.6500 114.9000 56.3500 115.6000 ;
      RECT 54.6500 114.9000 55.3500 115.6000 ;
      RECT 53.6500 114.9000 54.3500 115.6000 ;
      RECT 52.6500 114.9000 53.3500 115.6000 ;
      RECT 51.6500 114.9000 52.3500 115.6000 ;
      RECT 50.6500 114.9000 51.3500 115.6000 ;
      RECT 49.6500 114.9000 50.3500 115.6000 ;
      RECT 48.6500 114.9000 49.3500 115.6000 ;
      RECT 47.6500 114.9000 48.3500 115.6000 ;
      RECT 46.6500 114.9000 47.3500 115.6000 ;
      RECT 45.6500 114.9000 46.3500 115.6000 ;
      RECT 44.6500 114.9000 45.3500 115.6000 ;
      RECT 43.6500 114.9000 44.3500 115.6000 ;
      RECT 42.6500 114.9000 43.3500 115.6000 ;
      RECT 41.6500 114.9000 42.3500 115.6000 ;
      RECT 40.6500 114.9000 41.3500 115.6000 ;
      RECT 39.6500 114.9000 40.3500 115.6000 ;
      RECT 38.6500 114.9000 39.3500 115.6000 ;
      RECT 37.6500 114.9000 38.3500 115.6000 ;
      RECT 36.6500 114.9000 37.3500 115.6000 ;
      RECT 35.6500 114.9000 36.3500 115.6000 ;
      RECT 34.6500 114.9000 35.3500 115.6000 ;
      RECT 33.6500 114.9000 34.3500 115.6000 ;
      RECT 32.6500 114.9000 33.3500 115.6000 ;
      RECT 31.6500 114.9000 32.3500 115.6000 ;
      RECT 30.6500 114.9000 31.3500 115.6000 ;
      RECT 29.6500 114.9000 30.3500 115.6000 ;
      RECT 28.6500 114.9000 29.3500 115.6000 ;
      RECT 27.6500 114.9000 28.3500 115.6000 ;
      RECT 26.6500 114.9000 27.3500 115.6000 ;
      RECT 0.0000 114.9000 26.3500 115.6000 ;
      RECT 0.0000 0.7000 116.4000 114.9000 ;
      RECT 89.6500 0.0000 116.4000 0.7000 ;
      RECT 88.6500 0.0000 89.3500 0.7000 ;
      RECT 87.6500 0.0000 88.3500 0.7000 ;
      RECT 86.6500 0.0000 87.3500 0.7000 ;
      RECT 85.6500 0.0000 86.3500 0.7000 ;
      RECT 84.6500 0.0000 85.3500 0.7000 ;
      RECT 83.6500 0.0000 84.3500 0.7000 ;
      RECT 82.6500 0.0000 83.3500 0.7000 ;
      RECT 81.6500 0.0000 82.3500 0.7000 ;
      RECT 80.6500 0.0000 81.3500 0.7000 ;
      RECT 79.6500 0.0000 80.3500 0.7000 ;
      RECT 78.6500 0.0000 79.3500 0.7000 ;
      RECT 77.6500 0.0000 78.3500 0.7000 ;
      RECT 76.6500 0.0000 77.3500 0.7000 ;
      RECT 75.6500 0.0000 76.3500 0.7000 ;
      RECT 74.6500 0.0000 75.3500 0.7000 ;
      RECT 73.6500 0.0000 74.3500 0.7000 ;
      RECT 72.6500 0.0000 73.3500 0.7000 ;
      RECT 71.6500 0.0000 72.3500 0.7000 ;
      RECT 70.6500 0.0000 71.3500 0.7000 ;
      RECT 69.6500 0.0000 70.3500 0.7000 ;
      RECT 68.6500 0.0000 69.3500 0.7000 ;
      RECT 67.6500 0.0000 68.3500 0.7000 ;
      RECT 66.6500 0.0000 67.3500 0.7000 ;
      RECT 65.6500 0.0000 66.3500 0.7000 ;
      RECT 64.6500 0.0000 65.3500 0.7000 ;
      RECT 63.6500 0.0000 64.3500 0.7000 ;
      RECT 62.6500 0.0000 63.3500 0.7000 ;
      RECT 61.6500 0.0000 62.3500 0.7000 ;
      RECT 60.6500 0.0000 61.3500 0.7000 ;
      RECT 59.6500 0.0000 60.3500 0.7000 ;
      RECT 58.6500 0.0000 59.3500 0.7000 ;
      RECT 57.6500 0.0000 58.3500 0.7000 ;
      RECT 56.6500 0.0000 57.3500 0.7000 ;
      RECT 55.6500 0.0000 56.3500 0.7000 ;
      RECT 54.6500 0.0000 55.3500 0.7000 ;
      RECT 53.6500 0.0000 54.3500 0.7000 ;
      RECT 52.6500 0.0000 53.3500 0.7000 ;
      RECT 51.6500 0.0000 52.3500 0.7000 ;
      RECT 50.6500 0.0000 51.3500 0.7000 ;
      RECT 49.6500 0.0000 50.3500 0.7000 ;
      RECT 48.6500 0.0000 49.3500 0.7000 ;
      RECT 47.6500 0.0000 48.3500 0.7000 ;
      RECT 46.6500 0.0000 47.3500 0.7000 ;
      RECT 45.6500 0.0000 46.3500 0.7000 ;
      RECT 44.6500 0.0000 45.3500 0.7000 ;
      RECT 43.6500 0.0000 44.3500 0.7000 ;
      RECT 42.6500 0.0000 43.3500 0.7000 ;
      RECT 41.6500 0.0000 42.3500 0.7000 ;
      RECT 40.6500 0.0000 41.3500 0.7000 ;
      RECT 39.6500 0.0000 40.3500 0.7000 ;
      RECT 38.6500 0.0000 39.3500 0.7000 ;
      RECT 37.6500 0.0000 38.3500 0.7000 ;
      RECT 36.6500 0.0000 37.3500 0.7000 ;
      RECT 35.6500 0.0000 36.3500 0.7000 ;
      RECT 34.6500 0.0000 35.3500 0.7000 ;
      RECT 33.6500 0.0000 34.3500 0.7000 ;
      RECT 32.6500 0.0000 33.3500 0.7000 ;
      RECT 31.6500 0.0000 32.3500 0.7000 ;
      RECT 30.6500 0.0000 31.3500 0.7000 ;
      RECT 29.6500 0.0000 30.3500 0.7000 ;
      RECT 28.6500 0.0000 29.3500 0.7000 ;
      RECT 27.6500 0.0000 28.3500 0.7000 ;
      RECT 26.6500 0.0000 27.3500 0.7000 ;
      RECT 0.0000 0.0000 26.3500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 70.1500 116.4000 115.6000 ;
      RECT 0.7000 69.8500 116.4000 70.1500 ;
      RECT 0.0000 66.1500 116.4000 69.8500 ;
      RECT 0.7000 65.8500 116.4000 66.1500 ;
      RECT 0.0000 62.1500 116.4000 65.8500 ;
      RECT 0.7000 61.8500 116.4000 62.1500 ;
      RECT 0.0000 58.1500 116.4000 61.8500 ;
      RECT 0.7000 57.8500 116.4000 58.1500 ;
      RECT 0.0000 54.1500 116.4000 57.8500 ;
      RECT 0.7000 53.8500 116.4000 54.1500 ;
      RECT 0.0000 50.1500 116.4000 53.8500 ;
      RECT 0.7000 49.8500 116.4000 50.1500 ;
      RECT 0.0000 46.1500 116.4000 49.8500 ;
      RECT 0.7000 45.8500 116.4000 46.1500 ;
      RECT 0.0000 0.0000 116.4000 45.8500 ;
    LAYER M4 ;
      RECT 0.0000 114.2650 116.4000 115.6000 ;
      RECT 104.8200 114.1000 116.4000 114.2650 ;
      RECT 88.6000 114.1000 101.8200 114.2650 ;
      RECT 72.3800 114.1000 85.6000 114.2650 ;
      RECT 56.1600 114.1000 69.3800 114.2650 ;
      RECT 39.9400 114.1000 53.1600 114.2650 ;
      RECT 23.7200 114.1000 36.9400 114.2650 ;
      RECT 7.5000 114.1000 20.7200 114.2650 ;
      RECT 111.8200 1.5000 116.4000 114.1000 ;
      RECT 104.8200 1.5000 108.8200 114.1000 ;
      RECT 95.6000 1.5000 101.8200 114.1000 ;
      RECT 88.6000 1.5000 92.6000 114.1000 ;
      RECT 79.3800 1.5000 85.6000 114.1000 ;
      RECT 72.3800 1.5000 76.3800 114.1000 ;
      RECT 63.1600 1.5000 69.3800 114.1000 ;
      RECT 56.1600 1.5000 60.1600 114.1000 ;
      RECT 46.9400 1.5000 53.1600 114.1000 ;
      RECT 39.9400 1.5000 43.9400 114.1000 ;
      RECT 30.7200 1.5000 36.9400 114.1000 ;
      RECT 23.7200 1.5000 27.7200 114.1000 ;
      RECT 14.5000 1.5000 20.7200 114.1000 ;
      RECT 7.5000 1.5000 11.5000 114.1000 ;
      RECT 104.8200 1.3350 116.4000 1.5000 ;
      RECT 88.6000 1.3350 101.8200 1.5000 ;
      RECT 72.3800 1.3350 85.6000 1.5000 ;
      RECT 56.1600 1.3350 69.3800 1.5000 ;
      RECT 39.9400 1.3350 53.1600 1.5000 ;
      RECT 23.7200 1.3350 36.9400 1.5000 ;
      RECT 7.5000 1.3350 20.7200 1.5000 ;
      RECT 0.0000 1.3350 4.5000 114.2650 ;
      RECT 0.0000 0.0000 116.4000 1.3350 ;
  END
END sram_w8_64b

END LIBRARY
